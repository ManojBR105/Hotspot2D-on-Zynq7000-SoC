`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/02/2023 09:32:46 PM
// Design Name: 
// Module Name: Testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Testbench();

    parameter DATA_WIDTH = 32;

    reg                           aclk;
    reg                           axi_resetn;
    //temp data interface
    reg   [DATA_WIDTH-1:0]        s_axis_temp_data; //[c,n,s,e,w]
    wire                          s_axis_temp_ready;
    reg                           s_axis_temp_valid;
    
    //power data interface
    reg   [DATA_WIDTH-1:0]        s_axis_power_data;
    wire                          s_axis_power_ready;
    reg                           s_axis_power_valid;
    
    //result interface
    wire  [DATA_WIDTH*4-1:0]      m_axis_result_data;
    reg                           m_axis_result_ready;
    wire                          m_axis_result_valid;
    //config data
    reg   [DATA_WIDTH-1:0]        cns;
    reg   [DATA_WIDTH-1:0]        cwe;
    reg   [DATA_WIDTH-1:0]        cc;
    reg   [DATA_WIDTH-1:0]        Cap_1;
    reg   [DATA_WIDTH-1:0]        c_amb;
    
    reg    [DATA_WIDTH-1:0] temp_data[0:4999];
    reg    [DATA_WIDTH-1:0] power_data[0:4999];
    
    wire   [DATA_WIDTH*2-1:0]        out_temp;
    wire   [DATA_WIDTH*2-1:0]        out_power;
    wire   [DATA_WIDTH-1:0]        out_temp_32;
    
    wire   [DATA_WIDTH-1:0]        out_temp_fp;
        
    assign out_temp = m_axis_result_data[63:0];
    assign out_power = m_axis_result_data[95:64];
    assign out_temp_32 = out_temp[53:22];
    
    //testbench data store
    integer temp_counter;
    integer power_counter;
    
    wire ready_float_to_unit;
    wire valid_from_fp;
    
    sodaWithHotSpot #(.DATA_WIDTH(32),
                        .INT_WIDTH(10),
                        .FLOAT_WIDTH(22),
                        .SIZE(512)) sodaWithHotSpot_inst (
                        .aclk(aclk),
                        .axi_resetn(axi_resetn),
                        //temp data interface
                        .s_axis_temp_data(s_axis_temp_data), 
                        .s_axis_temp_ready(s_axis_temp_ready),
                        .s_axis_temp_valid(s_axis_temp_valid),
                        //power data interface
                        .s_axis_power_data(s_axis_power_data),
                        .s_axis_power_ready(s_axis_power_ready),
                        .s_axis_power_valid(s_axis_power_valid),
                        //output temp interface
                        .m_axis_result_data(m_axis_result_data), //{power,temp}
                        .m_axis_result_ready(ready_float_to_unit),
                        .m_axis_result_valid(m_axis_result_valid),
                        //config data
                        .cns(cns),
                        .cwe(cwe),
                        .cc(cc),
                        .Cap_1(Cap_1),
                        .c_amb(c_amb) 

    );
    
    floating_point_0 your_instance_name (
      .aclk(aclk),                                  // input wire aclk
      .s_axis_a_tvalid(m_axis_result_valid),            // input wire s_axis_a_tvalid
      .s_axis_a_tready(ready_float_to_unit),            // output wire s_axis_a_tready
      .s_axis_a_tdata(out_temp),              // input wire [63 : 0] s_axis_a_tdata
      .m_axis_result_tvalid(valid_from_fp),  // output wire m_axis_result_tvalid
      .m_axis_result_tready(m_axis_result_ready),  // input wire m_axis_result_tready
      .m_axis_result_tdata(out_temp_fp)    // output wire [31 : 0] m_axis_result_tdata
    );
    
    initial begin
        /*temp_data[0] = 32'h01c00000; //7
        temp_data[1] = 32'h02000000; //8
        temp_data[2] = 32'h02400000; //9
        temp_data[3] = 32'h02800000; //10
        temp_data[4] = 32'h02c00000; //11
        temp_data[5] = 32'h06c00000; //27
        temp_data[6] = 32'h07c00000; //31
        temp_data[7] = 32'h04c00000; //19
        temp_data[8] = 32'h05400000; //21
        temp_data[9] = 32'h04400000; //17
        
        
        power_data[0] = 32'h03000000;
        power_data[1] = 32'h09000000;
        power_data[2] = 32'h04cccccd;
        power_data[3] = 32'h02c00000;
        power_data[4] = 32'h030f11b6;
        power_data[5] = 32'h0096b4d0;
        power_data[6] = 32'h04cf1206;
        power_data[7] = 32'h03d7aa8b;
        power_data[8] = 32'h031700a8;
        power_data[9] = 32'h05ecb2c8;  
        */
        
        temp_counter = 0;     
        power_counter = 0;
    end
    
    //clock handle
    initial begin
        aclk = 0;
        forever #2 aclk = ~aclk;
    end
    
    //reset handle
    initial begin
        axi_resetn = 0;
        #7;
        axi_resetn = 1;
    end
    
    //passing temp data
    always @(negedge aclk) begin
        if(~axi_resetn) begin
            s_axis_temp_data <= {DATA_WIDTH{1'b0}};
        end
        else begin
            if(s_axis_temp_ready & s_axis_temp_valid) begin
                s_axis_temp_data <= temp_data[temp_counter];
                if(temp_counter == 512*512+512) 
                    temp_counter = 0;
                else
                    temp_counter=temp_counter+1;
            end
        end
    end
    
    
    //passing power data
    always @(negedge aclk) begin
        if(~axi_resetn) begin
            s_axis_power_data <= {DATA_WIDTH*{1'b0}};
        end
        else begin
            if(s_axis_power_ready & s_axis_power_valid) begin
                s_axis_power_data <= power_data[power_counter];
                if(power_counter == 512*512+512) 
                    power_counter = 0;
                else
                    power_counter=power_counter+1;
            end
        end
    end
    
    //control validity of temp data
    initial begin
        s_axis_temp_valid = 0;
        #24;
        s_axis_temp_valid = 1;
        s_axis_temp_data <= temp_data[0];
        #16;
        s_axis_temp_valid = 0;
        #8;
        s_axis_temp_valid = 1;
        #20;
        s_axis_temp_valid = 0;
        #8;
        s_axis_temp_valid = 1;
        #20;
        s_axis_temp_valid = 0;
        #8;
        s_axis_temp_valid = 1;
        #68;
        s_axis_temp_valid = 0;
        #68;
        s_axis_temp_valid = 1;
    end
    
    //control validity of power data
    initial begin
        s_axis_power_valid = 0;
        #12;
        s_axis_power_valid = 1;
        s_axis_power_data <= power_data[0];
        #20;
        s_axis_power_valid = 0;
        #8;
        s_axis_power_valid = 1;
        #20;
        s_axis_power_valid = 0;
        #8;
        s_axis_power_valid = 1;
        #20;
        s_axis_power_valid = 0;
        #8;
        s_axis_power_valid = 1;
        #68;
        s_axis_power_valid = 0;
        #68;
        s_axis_power_valid = 1;
    end
    
    
    //handling master ready
    initial begin
        m_axis_result_ready = 0;
        #7;
        m_axis_result_ready = 1;
        #24;
        m_axis_result_ready = 0;
        #12;
        m_axis_result_ready = 1;
        #4;
        m_axis_result_ready = 0;
        #16;
        m_axis_result_ready = 1;
        #48;
        m_axis_result_ready = 0;
        #16;
        m_axis_result_ready = 1;
        
    end
    
    //config handle
    initial begin
        cns = 32'h00000596; //0.125
        cwe = 32'h00000596; //0.256
        cc = 32'h003fe99f; //0.856
        Cap_1 = 32'h000037eb; //1.864
        c_amb = 32'h0000022e; //82.94
    end
   
    //simulation time handle
    initial begin
        #4000000000;
        $finish;
    end
    

    initial begin
temp_data[0] = 32'h50f71bdf;
temp_data[1] = 32'h50f72820;
temp_data[2] = 32'h50f73f70;
temp_data[3] = 32'h50f7609a;
temp_data[4] = 32'h50f78a8f;
temp_data[5] = 32'h50f7bc51;
temp_data[6] = 32'h50f7f50a;
temp_data[7] = 32'h50f833f4;
temp_data[8] = 32'h50f87860;
temp_data[9] = 32'h50f8c1a9;
temp_data[10] = 32'h50f90f45;
temp_data[11] = 32'h50f960b7;
temp_data[12] = 32'h50f9b58d;
temp_data[13] = 32'h50fa0d5f;
temp_data[14] = 32'h50fa67d3;
temp_data[15] = 32'h50fac497;
temp_data[16] = 32'h50fb2364;
temp_data[17] = 32'h50fb83f9;
temp_data[18] = 32'h50fbe61d;
temp_data[19] = 32'h50fc499d;
temp_data[20] = 32'h50fcae47;
temp_data[21] = 32'h50fd13f5;
temp_data[22] = 32'h50fd7a85;
temp_data[23] = 32'h50fde1d6;
temp_data[24] = 32'h50fe49cb;
temp_data[25] = 32'h50feb24a;
temp_data[26] = 32'h50ff1b3f;
temp_data[27] = 32'h50ff8499;
temp_data[28] = 32'h50ffee42;
temp_data[29] = 32'h5100582e;
temp_data[30] = 32'h5100c250;
temp_data[31] = 32'h51012c9d;
temp_data[32] = 32'h5101970b;
temp_data[33] = 32'h51020197;
temp_data[34] = 32'h51026c33;
temp_data[35] = 32'h5102d6e0;
temp_data[36] = 32'h51034196;
temp_data[37] = 32'h5103ac4f;
temp_data[38] = 32'h5104170d;
temp_data[39] = 32'h510481cb;
temp_data[40] = 32'h5104ec85;
temp_data[41] = 32'h51055743;
temp_data[42] = 32'h5105c1fd;
temp_data[43] = 32'h51062cb6;
temp_data[44] = 32'h51069770;
temp_data[45] = 32'h51070225;
temp_data[46] = 32'h51076cdf;
temp_data[47] = 32'h5107d79d;
temp_data[48] = 32'h5108425f;
temp_data[49] = 32'h5108ad2a;
temp_data[50] = 32'h510917fc;
temp_data[51] = 32'h510982dc;
temp_data[52] = 32'h5109edcc;
temp_data[53] = 32'h510a58c9;
temp_data[54] = 32'h510ac3df;
temp_data[55] = 32'h510b2f0e;
temp_data[56] = 32'h510b9a56;
temp_data[57] = 32'h510c05c0;
temp_data[58] = 32'h510c714c;
temp_data[59] = 32'h510cdd01;
temp_data[60] = 32'h510d48dc;
temp_data[61] = 32'h510db4ea;
temp_data[62] = 32'h510e2125;
temp_data[63] = 32'h510e8d9b;
temp_data[64] = 32'h510efa48;
temp_data[65] = 32'h510f6734;
temp_data[66] = 32'h510fd467;
temp_data[67] = 32'h511041dd;
temp_data[68] = 32'h5110afa3;
temp_data[69] = 32'h51111db8;
temp_data[70] = 32'h51118c22;
temp_data[71] = 32'h5111fae3;
temp_data[72] = 32'h51126a05;
temp_data[73] = 32'h5112d98c;
temp_data[74] = 32'h51134977;
temp_data[75] = 32'h5113b9d4;
temp_data[76] = 32'h51142aa2;
temp_data[77] = 32'h51149be9;
temp_data[78] = 32'h51150daa;
temp_data[79] = 32'h51157ff1;
temp_data[80] = 32'h5115f2bf;
temp_data[81] = 32'h5116661b;
temp_data[82] = 32'h5116da0a;
temp_data[83] = 32'h51174e94;
temp_data[84] = 32'h5117c3bd;
temp_data[85] = 32'h5118398a;
temp_data[86] = 32'h5118b008;
temp_data[87] = 32'h51192739;
temp_data[88] = 32'h51199f1f;
temp_data[89] = 32'h511a17ca;
temp_data[90] = 32'h511a913f;
temp_data[91] = 32'h511b0b80;
temp_data[92] = 32'h511b869c;
temp_data[93] = 32'h511c0297;
temp_data[94] = 32'h511c7f78;
temp_data[95] = 32'h511cfd48;
temp_data[96] = 32'h511d7c13;
temp_data[97] = 32'h511dfbdf;
temp_data[98] = 32'h511e7cb7;
temp_data[99] = 32'h511efea4;
temp_data[100] = 32'h511f81b2;
temp_data[101] = 32'h512005ea;
temp_data[102] = 32'h51208b59;
temp_data[103] = 32'h51211206;
temp_data[104] = 32'h51219a02;
temp_data[105] = 32'h51222357;
temp_data[106] = 32'h5122ae14;
temp_data[107] = 32'h51233a4b;
temp_data[108] = 32'h5123c800;
temp_data[109] = 32'h51245747;
temp_data[110] = 32'h5124e836;
temp_data[111] = 32'h51257ad1;
temp_data[112] = 32'h51260f34;
temp_data[113] = 32'h5126a56e;
temp_data[114] = 32'h51273d92;
temp_data[115] = 32'h5127d7ae;
temp_data[116] = 32'h512873de;
temp_data[117] = 32'h51291238;
temp_data[118] = 32'h5129b2cc;
temp_data[119] = 32'h512a55b4;
temp_data[120] = 32'h512afb0d;
temp_data[121] = 32'h512ba2e8;
temp_data[122] = 32'h512c4d62;
temp_data[123] = 32'h512cfa98;
temp_data[124] = 32'h512daaa4;
temp_data[125] = 32'h512e5da2;
temp_data[126] = 32'h512f13ad;
temp_data[127] = 32'h512fcce6;
temp_data[128] = 32'h51308965;
temp_data[129] = 32'h51314949;
temp_data[130] = 32'h51320cae;
temp_data[131] = 32'h5132d3b7;
temp_data[132] = 32'h51339e73;
temp_data[133] = 32'h51346d05;
temp_data[134] = 32'h51353f85;
temp_data[135] = 32'h51361605;
temp_data[136] = 32'h5136f095;
temp_data[137] = 32'h5137cf4a;
temp_data[138] = 32'h5138b229;
temp_data[139] = 32'h51399939;
temp_data[140] = 32'h513a8477;
temp_data[141] = 32'h513b73d6;
temp_data[142] = 32'h513c6745;
temp_data[143] = 32'h513d5eab;
temp_data[144] = 32'h513e59e2;
temp_data[145] = 32'h513f58b0;
temp_data[146] = 32'h51405ad9;
temp_data[147] = 32'h5141600f;
temp_data[148] = 32'h514267f5;
temp_data[149] = 32'h51437222;
temp_data[150] = 32'h51447e17;
temp_data[151] = 32'h51458b48;
temp_data[152] = 32'h51469918;
temp_data[153] = 32'h5147a6df;
temp_data[154] = 32'h5148b3e1;
temp_data[155] = 32'h5149bf59;
temp_data[156] = 32'h514ac871;
temp_data[157] = 32'h514bcfe1;
temp_data[158] = 32'h514cdb40;
temp_data[159] = 32'h514de9af;
temp_data[160] = 32'h514efa66;
temp_data[161] = 32'h51500ca2;
temp_data[162] = 32'h51511fb4;
temp_data[163] = 32'h51523305;
temp_data[164] = 32'h51534602;
temp_data[165] = 32'h51545832;
temp_data[166] = 32'h5155692b;
temp_data[167] = 32'h51567892;
temp_data[168] = 32'h51578627;
temp_data[169] = 32'h515891b0;
temp_data[170] = 32'h51599b02;
temp_data[171] = 32'h515aa20a;
temp_data[172] = 32'h515ba6bd;
temp_data[173] = 32'h515ca922;
temp_data[174] = 32'h515da93f;
temp_data[175] = 32'h515ea737;
temp_data[176] = 32'h515fa32f;
temp_data[177] = 32'h51609d56;
temp_data[178] = 32'h516195e1;
temp_data[179] = 32'h51628d19;
temp_data[180] = 32'h51638345;
temp_data[181] = 32'h516478b8;
temp_data[182] = 32'h51656dd2;
temp_data[183] = 32'h516662f6;
temp_data[184] = 32'h5167588e;
temp_data[185] = 32'h51684f16;
temp_data[186] = 32'h5169470f;
temp_data[187] = 32'h516a40ff;
temp_data[188] = 32'h516b3d81;
temp_data[189] = 32'h516c3d3a;
temp_data[190] = 32'h516d40d9;
temp_data[191] = 32'h516e491f;
temp_data[192] = 32'h516f56de;
temp_data[193] = 32'h51706af4;
temp_data[194] = 32'h51718662;
temp_data[195] = 32'h5172aa2e;
temp_data[196] = 32'h5173d784;
temp_data[197] = 32'h51750fae;
temp_data[198] = 32'h51765409;
temp_data[199] = 32'h5177a61e;
temp_data[200] = 32'h5179079e;
temp_data[201] = 32'h517a7a63;
temp_data[202] = 32'h517c007a;
temp_data[203] = 32'h517d9c24;
temp_data[204] = 32'h517f4fdf;
temp_data[205] = 32'h51811e6d;
temp_data[206] = 32'h51830ad9;
temp_data[207] = 32'h5185187e;
temp_data[208] = 32'h51874b1f;
temp_data[209] = 32'h5189a6d7;
temp_data[210] = 32'h518c3040;
temp_data[211] = 32'h518eec63;
temp_data[212] = 32'h5191e0df;
temp_data[213] = 32'h519513ec;
temp_data[214] = 32'h51988c6d;
temp_data[215] = 32'h519c5200;
temp_data[216] = 32'h51a06d1a;
temp_data[217] = 32'h51a4e70c;
temp_data[218] = 32'h51a9ca32;
temp_data[219] = 32'h51af21fb;
temp_data[220] = 32'h51b4fb0d;
temp_data[221] = 32'h51bb6367;
temp_data[222] = 32'h51c26a7b;
temp_data[223] = 32'h51ca215c;
temp_data[224] = 32'h51d29ae5;
temp_data[225] = 32'h51dbebea;
temp_data[226] = 32'h51e62b67;
temp_data[227] = 32'h51f172da;
temp_data[228] = 32'h51fc074f;
temp_data[229] = 32'h52058d58;
temp_data[230] = 32'h520e1c76;
temp_data[231] = 32'h5215c99f;
temp_data[232] = 32'h521ca783;
temp_data[233] = 32'h5222c6b0;
temp_data[234] = 32'h522835b9;
temp_data[235] = 32'h522d0165;
temp_data[236] = 32'h523134ca;
temp_data[237] = 32'h5234d95e;
temp_data[238] = 32'h5237f723;
temp_data[239] = 32'h523a94a7;
temp_data[240] = 32'h523cb720;
temp_data[241] = 32'h523e6278;
temp_data[242] = 32'h523f995f;
temp_data[243] = 32'h52405d3a;
temp_data[244] = 32'h5240ae47;
temp_data[245] = 32'h52408b8b;
temp_data[246] = 32'h523ff2d0;
temp_data[247] = 32'h523ee0b1;
temp_data[248] = 32'h523d507a;
temp_data[249] = 32'h523b3c36;
temp_data[250] = 32'h52389c8d;
temp_data[251] = 32'h523568b6;
temp_data[252] = 32'h52319668;
temp_data[253] = 32'h522d19c6;
temp_data[254] = 32'h5227e52a;
temp_data[255] = 32'h5221e914;
temp_data[256] = 32'h521b13e8;
temp_data[257] = 32'h5215276b;
temp_data[258] = 32'h52101223;
temp_data[259] = 32'h520bc4b9;
temp_data[260] = 32'h520831d7;
temp_data[261] = 32'h52054e01;
temp_data[262] = 32'h52030f6f;
temp_data[263] = 32'h52016dfc;
temp_data[264] = 32'h5200630b;
temp_data[265] = 32'h51ffe97d;
temp_data[266] = 32'h51fffda0;
temp_data[267] = 32'h52009d34;
temp_data[268] = 32'h5201c754;
temp_data[269] = 32'h52037c78;
temp_data[270] = 32'h5205be8c;
temp_data[271] = 32'h520890da;
temp_data[272] = 32'h520bf82f;
temp_data[273] = 32'h520ffad3;
temp_data[274] = 32'h5214a0ae;
temp_data[275] = 32'h5219f34d;
temp_data[276] = 32'h521ffe15;
temp_data[277] = 32'h5226ce46;
temp_data[278] = 32'h522e7336;
temp_data[279] = 32'h5236fe7a;
temp_data[280] = 32'h5240840e;
temp_data[281] = 32'h524b1a87;
temp_data[282] = 32'h5256db6a;
temp_data[283] = 32'h5263e350;
temp_data[284] = 32'h52725254;
temp_data[285] = 32'h52824c51;
temp_data[286] = 32'h5293f944;
temp_data[287] = 32'h52a785ba;
temp_data[288] = 32'h52bd2353;
temp_data[289] = 32'h52d5091c;
temp_data[290] = 32'h52ef7443;
temp_data[291] = 32'h530ca89c;
temp_data[292] = 32'h532cf156;
temp_data[293] = 32'h5350a1b6;
temp_data[294] = 32'h537815df;
temp_data[295] = 32'h53a3b3cc;
temp_data[296] = 32'h53d3ec39;
temp_data[297] = 32'h54093c15;
temp_data[298] = 32'h543f99d0;
temp_data[299] = 32'h5470b4ab;
temp_data[300] = 32'h549d0c28;
temp_data[301] = 32'h54c5134d;
temp_data[302] = 32'h54e93205;
temp_data[303] = 32'h5509c64c;
temp_data[304] = 32'h552724f2;
temp_data[305] = 32'h55419a91;
temp_data[306] = 32'h55596c3c;
temp_data[307] = 32'h556ed830;
temp_data[308] = 32'h55821676;
temp_data[309] = 32'h55935971;
temp_data[310] = 32'h55a2ce57;
temp_data[311] = 32'h55b09dbb;
temp_data[312] = 32'h55bcebe6;
temp_data[313] = 32'h55c7d93c;
temp_data[314] = 32'h55d18290;
temp_data[315] = 32'h55da0179;
temp_data[316] = 32'h55e16c94;
temp_data[317] = 32'h55e7d7ba;
temp_data[318] = 32'h55ed5443;
temp_data[319] = 32'h55f1f12c;
temp_data[320] = 32'h55f5bb45;
temp_data[321] = 32'h55f8bd55;
temp_data[322] = 32'h55fb003b;
temp_data[323] = 32'h55fc8af8;
temp_data[324] = 32'h55fd62d4;
temp_data[325] = 32'h55fd8b6e;
temp_data[326] = 32'h55fd06b3;
temp_data[327] = 32'h55fbd4f6;
temp_data[328] = 32'h55f9f4e8;
temp_data[329] = 32'h55f76399;
temp_data[330] = 32'h55f41c76;
temp_data[331] = 32'h55f01922;
temp_data[332] = 32'h55eb518b;
temp_data[333] = 32'h55e5bbb6;
temp_data[334] = 32'h55df4ba9;
temp_data[335] = 32'h55d7f35a;
temp_data[336] = 32'h55cfa26e;
temp_data[337] = 32'h55c64628;
temp_data[338] = 32'h55bbc921;
temp_data[339] = 32'h55b01316;
temp_data[340] = 32'h55a308a2;
temp_data[341] = 32'h55948af8;
temp_data[342] = 32'h5584778e;
temp_data[343] = 32'h5572a7c6;
temp_data[344] = 32'h555ef080;
temp_data[345] = 32'h554921ab;
temp_data[346] = 32'h553105cd;
temp_data[347] = 32'h55166174;
temp_data[348] = 32'h54f8f29d;
temp_data[349] = 32'h54d8700d;
temp_data[350] = 32'h54b4889c;
temp_data[351] = 32'h548ce25d;
temp_data[352] = 32'h546119ce;
temp_data[353] = 32'h5430c0ca;
temp_data[354] = 32'h53fb5d79;
temp_data[355] = 32'h53c068a9;
temp_data[356] = 32'h5388cd92;
temp_data[357] = 32'h53565f78;
temp_data[358] = 32'h53289f45;
temp_data[359] = 32'h52ff19fc;
temp_data[360] = 32'h52d967ae;
temp_data[361] = 32'h52b72a41;
temp_data[362] = 32'h52980c9e;
temp_data[363] = 32'h527bc1ce;
temp_data[364] = 32'h5262044b;
temp_data[365] = 32'h524a9531;
temp_data[366] = 32'h52353bbc;
temp_data[367] = 32'h5221c4a0;
temp_data[368] = 32'h5210018a;
temp_data[369] = 32'h51ffc8b4;
temp_data[370] = 32'h51f0f45e;
temp_data[371] = 32'h51e3627c;
temp_data[372] = 32'h51d6f45e;
temp_data[373] = 32'h51cb8e47;
temp_data[374] = 32'h51c1173c;
temp_data[375] = 32'h51b778b3;
temp_data[376] = 32'h51ae9e52;
temp_data[377] = 32'h51a675c9;
temp_data[378] = 32'h519eee80;
temp_data[379] = 32'h5197f994;
temp_data[380] = 32'h51918987;
temp_data[381] = 32'h518b9232;
temp_data[382] = 32'h5186089a;
temp_data[383] = 32'h5180e2d6;
temp_data[384] = 32'h517c17f0;
temp_data[385] = 32'h51779fd3;
temp_data[386] = 32'h51737336;
temp_data[387] = 32'h516f8b76;
temp_data[388] = 32'h516be29b;
temp_data[389] = 32'h5168733f;
temp_data[390] = 32'h5165387e;
temp_data[391] = 32'h51622de4;
temp_data[392] = 32'h515f4f76;
temp_data[393] = 32'h515c9985;
temp_data[394] = 32'h515a08d1;
temp_data[395] = 32'h51579a4e;
temp_data[396] = 32'h51554b4d;
temp_data[397] = 32'h51531950;
temp_data[398] = 32'h51510219;
temp_data[399] = 32'h514f039f;
temp_data[400] = 32'h514d1c00;
temp_data[401] = 32'h514b4990;
temp_data[402] = 32'h51498ac2;
temp_data[403] = 32'h5147de27;
temp_data[404] = 32'h5146427c;
temp_data[405] = 32'h5144b68d;
temp_data[406] = 32'h5143394b;
temp_data[407] = 32'h5141c9b4;
temp_data[408] = 32'h514066e8;
temp_data[409] = 32'h513f100a;
temp_data[410] = 32'h513dc459;
temp_data[411] = 32'h513c8327;
temp_data[412] = 32'h513b4bc7;
temp_data[413] = 32'h513a1da3;
temp_data[414] = 32'h5138f834;
temp_data[415] = 32'h5137daec;
temp_data[416] = 32'h5136c561;
temp_data[417] = 32'h5135b71c;
temp_data[418] = 32'h5134afb4;
temp_data[419] = 32'h5133aed1;
temp_data[420] = 32'h5132b414;
temp_data[421] = 32'h5131bf2b;
temp_data[422] = 32'h5130cfcc;
temp_data[423] = 32'h512fe5ac;
temp_data[424] = 32'h512f008a;
temp_data[425] = 32'h512e2029;
temp_data[426] = 32'h512d444e;
temp_data[427] = 32'h512c6cbe;
temp_data[428] = 32'h512b9946;
temp_data[429] = 32'h512ac9b8;
temp_data[430] = 32'h5129fde7;
temp_data[431] = 32'h512935a8;
temp_data[432] = 32'h512870d2;
temp_data[433] = 32'h5127af3a;
temp_data[434] = 32'h5126f0c3;
temp_data[435] = 32'h51263544;
temp_data[436] = 32'h51257ca2;
temp_data[437] = 32'h5124c6bd;
temp_data[438] = 32'h51241377;
temp_data[439] = 32'h512362b2;
temp_data[440] = 32'h5122b457;
temp_data[441] = 32'h5122084f;
temp_data[442] = 32'h51215e78;
temp_data[443] = 32'h5120b6c8;
temp_data[444] = 32'h5120111f;
temp_data[445] = 32'h511f6d6e;
temp_data[446] = 32'h511ecb9b;
temp_data[447] = 32'h511e2b99;
temp_data[448] = 32'h511d8d54;
temp_data[449] = 32'h511cf0bb;
temp_data[450] = 32'h511c55b9;
temp_data[451] = 32'h511bbc41;
temp_data[452] = 32'h511b2442;
temp_data[453] = 32'h511a8db0;
temp_data[454] = 32'h5119f87b;
temp_data[455] = 32'h51196499;
temp_data[456] = 32'h5118d1f6;
temp_data[457] = 32'h51184085;
temp_data[458] = 32'h5117b042;
temp_data[459] = 32'h5117211d;
temp_data[460] = 32'h5116930c;
temp_data[461] = 32'h51160603;
temp_data[462] = 32'h511579f6;
temp_data[463] = 32'h5114eee1;
temp_data[464] = 32'h511464bb;
temp_data[465] = 32'h5113db73;
temp_data[466] = 32'h5113530d;
temp_data[467] = 32'h5112cb79;
temp_data[468] = 32'h511244b3;
temp_data[469] = 32'h5111beb6;
temp_data[470] = 32'h5111397a;
temp_data[471] = 32'h5110b4fa;
temp_data[472] = 32'h51103138;
temp_data[473] = 32'h510fae29;
temp_data[474] = 32'h510f2bd0;
temp_data[475] = 32'h510eaa26;
temp_data[476] = 32'h510e2930;
temp_data[477] = 32'h510da8eb;
temp_data[478] = 32'h510d2956;
temp_data[479] = 32'h510caa7a;
temp_data[480] = 32'h510c2c56;
temp_data[481] = 32'h510baef3;
temp_data[482] = 32'h510b3255;
temp_data[483] = 32'h510ab689;
temp_data[484] = 32'h510a3b92;
temp_data[485] = 32'h5109c183;
temp_data[486] = 32'h5109486b;
temp_data[487] = 32'h5108d05b;
temp_data[488] = 32'h51085968;
temp_data[489] = 32'h5107e3a8;
temp_data[490] = 32'h51076f3b;
temp_data[491] = 32'h5106fc3b;
temp_data[492] = 32'h51068ad2;
temp_data[493] = 32'h51061b26;
temp_data[494] = 32'h5105ad60;
temp_data[495] = 32'h510541bc;
temp_data[496] = 32'h5104d86f;
temp_data[497] = 32'h510471bd;
temp_data[498] = 32'h51040ded;
temp_data[499] = 32'h5103ad58;
temp_data[500] = 32'h51035059;
temp_data[501] = 32'h5102f751;
temp_data[502] = 32'h5102a2be;
temp_data[503] = 32'h5102531e;
temp_data[504] = 32'h510208ff;
temp_data[505] = 32'h5101c509;
temp_data[506] = 32'h510187ec;
temp_data[507] = 32'h51015276;
temp_data[508] = 32'h51012581;
temp_data[509] = 32'h51010210;
temp_data[510] = 32'h5100e936;
temp_data[511] = 32'h5100dc27;
temp_data[512] = 32'h50f71961;
temp_data[513] = 32'h50f725a7;
temp_data[514] = 32'h50f73cfb;
temp_data[515] = 32'h50f75e2d;
temp_data[516] = 32'h50f78827;
temp_data[517] = 32'h50f7b9f1;
temp_data[518] = 32'h50f7f2b6;
temp_data[519] = 32'h50f831ad;
temp_data[520] = 32'h50f87621;
temp_data[521] = 32'h50f8bf7b;
temp_data[522] = 32'h50f90d24;
temp_data[523] = 32'h50f95ea6;
temp_data[524] = 32'h50f9b389;
temp_data[525] = 32'h50fa0b6b;
temp_data[526] = 32'h50fa65f1;
temp_data[527] = 32'h50fac2c6;
temp_data[528] = 32'h50fb21a3;
temp_data[529] = 32'h50fb824d;
temp_data[530] = 32'h50fbe482;
temp_data[531] = 32'h50fc480f;
temp_data[532] = 32'h50fcaccd;
temp_data[533] = 32'h50fd1290;
temp_data[534] = 32'h50fd7931;
temp_data[535] = 32'h50fde098;
temp_data[536] = 32'h50fe489d;
temp_data[537] = 32'h50feb131;
temp_data[538] = 32'h50ff1a3b;
temp_data[539] = 32'h50ff83a5;
temp_data[540] = 32'h50ffed63;
temp_data[541] = 32'h51005760;
temp_data[542] = 32'h5100c198;
temp_data[543] = 32'h51012bfa;
temp_data[544] = 32'h51019681;
temp_data[545] = 32'h5102011d;
temp_data[546] = 32'h51026bcf;
temp_data[547] = 32'h5102d691;
temp_data[548] = 32'h51034157;
temp_data[549] = 32'h5103ac2a;
temp_data[550] = 32'h510416f8;
temp_data[551] = 32'h510481cb;
temp_data[552] = 32'h5104ec9e;
temp_data[553] = 32'h51055771;
temp_data[554] = 32'h5105c240;
temp_data[555] = 32'h51062d0e;
temp_data[556] = 32'h510697dd;
temp_data[557] = 32'h510702ac;
temp_data[558] = 32'h51076d7a;
temp_data[559] = 32'h5107d84d;
temp_data[560] = 32'h51084324;
temp_data[561] = 32'h5108ae04;
temp_data[562] = 32'h510918ec;
temp_data[563] = 32'h510983e4;
temp_data[564] = 32'h5109eee5;
temp_data[565] = 32'h510a59fb;
temp_data[566] = 32'h510ac52a;
temp_data[567] = 32'h510b306e;
temp_data[568] = 32'h510b9bcc;
temp_data[569] = 32'h510c074f;
temp_data[570] = 32'h510c72ef;
temp_data[571] = 32'h510cdeb9;
temp_data[572] = 32'h510d4aae;
temp_data[573] = 32'h510db6d0;
temp_data[574] = 32'h510e2325;
temp_data[575] = 32'h510e8fb0;
temp_data[576] = 32'h510efc76;
temp_data[577] = 32'h510f697b;
temp_data[578] = 32'h510fd6c3;
temp_data[579] = 32'h51104452;
temp_data[580] = 32'h5110b22d;
temp_data[581] = 32'h51112058;
temp_data[582] = 32'h51118eda;
temp_data[583] = 32'h5111fdb5;
temp_data[584] = 32'h51126cf0;
temp_data[585] = 32'h5112dc90;
temp_data[586] = 32'h51134c94;
temp_data[587] = 32'h5113bd0a;
temp_data[588] = 32'h51142df1;
temp_data[589] = 32'h51149f4d;
temp_data[590] = 32'h5115112c;
temp_data[591] = 32'h51158388;
temp_data[592] = 32'h5115f66f;
temp_data[593] = 32'h511669e8;
temp_data[594] = 32'h5116ddf0;
temp_data[595] = 32'h51175293;
temp_data[596] = 32'h5117c7d6;
temp_data[597] = 32'h51183dc0;
temp_data[598] = 32'h5118b45b;
temp_data[599] = 32'h51192ba1;
temp_data[600] = 32'h5119a3a9;
temp_data[601] = 32'h511a1c6d;
temp_data[602] = 32'h511a95ff;
temp_data[603] = 32'h511b105e;
temp_data[604] = 32'h511b8b93;
temp_data[605] = 32'h511c07ab;
temp_data[606] = 32'h511c84a9;
temp_data[607] = 32'h511d0297;
temp_data[608] = 32'h511d8180;
temp_data[609] = 32'h511e016d;
temp_data[610] = 32'h511e8262;
temp_data[611] = 32'h511f0471;
temp_data[612] = 32'h511f879c;
temp_data[613] = 32'h51200bf6;
temp_data[614] = 32'h51209186;
temp_data[615] = 32'h51211855;
temp_data[616] = 32'h5121a073;
temp_data[617] = 32'h512229ed;
temp_data[618] = 32'h5122b4d0;
temp_data[619] = 32'h51234129;
temp_data[620] = 32'h5123cf03;
temp_data[621] = 32'h51245e74;
temp_data[622] = 32'h5124ef85;
temp_data[623] = 32'h5125824d;
temp_data[624] = 32'h512616d7;
temp_data[625] = 32'h5126ad3f;
temp_data[626] = 32'h5127458d;
temp_data[627] = 32'h5127dfdb;
temp_data[628] = 32'h51287c39;
temp_data[629] = 32'h51291ac1;
temp_data[630] = 32'h5129bb8c;
temp_data[631] = 32'h512a5eab;
temp_data[632] = 32'h512b043a;
temp_data[633] = 32'h512bac4f;
temp_data[634] = 32'h512c5708;
temp_data[635] = 32'h512d0481;
temp_data[636] = 32'h512db4d0;
temp_data[637] = 32'h512e6816;
temp_data[638] = 32'h512f1e71;
temp_data[639] = 32'h512fd7f9;
temp_data[640] = 32'h513094d1;
temp_data[641] = 32'h51315511;
temp_data[642] = 32'h513218db;
temp_data[643] = 32'h5132e04c;
temp_data[644] = 32'h5133ab7e;
temp_data[645] = 32'h51347a8d;
temp_data[646] = 32'h51354d90;
temp_data[647] = 32'h5136249e;
temp_data[648] = 32'h5136ffc9;
temp_data[649] = 32'h5137df26;
temp_data[650] = 32'h5138c2b9;
temp_data[651] = 32'h5139aa8b;
temp_data[652] = 32'h513a9696;
temp_data[653] = 32'h513b86d7;
temp_data[654] = 32'h513c7b3e;
temp_data[655] = 32'h513d73a8;
temp_data[656] = 32'h513e6ff4;
temp_data[657] = 32'h513f6fef;
temp_data[658] = 32'h51407358;
temp_data[659] = 32'h514179e6;
temp_data[660] = 32'h51428334;
temp_data[661] = 32'h51438ede;
temp_data[662] = 32'h51449c63;
temp_data[663] = 32'h5145ab32;
temp_data[664] = 32'h5146bab2;
temp_data[665] = 32'h5147ca3a;
temp_data[666] = 32'h5148d902;
temp_data[667] = 32'h5149e64b;
temp_data[668] = 32'h514af135;
temp_data[669] = 32'h514bfa7b;
temp_data[670] = 32'h514d07ab;
temp_data[671] = 32'h514e17e7;
temp_data[672] = 32'h514f2a5e;
temp_data[673] = 32'h51503e53;
temp_data[674] = 32'h51515311;
temp_data[675] = 32'h515267f9;
temp_data[676] = 32'h51537c7c;
temp_data[677] = 32'h5154901d;
temp_data[678] = 32'h5155a277;
temp_data[679] = 32'h5156b329;
temp_data[680] = 32'h5157c1f4;
temp_data[681] = 32'h5158ce9a;
temp_data[682] = 32'h5159d8f9;
temp_data[683] = 32'h515ae0fc;
temp_data[684] = 32'h515be697;
temp_data[685] = 32'h515ce9d1;
temp_data[686] = 32'h515deab3;
temp_data[687] = 32'h515ee964;
temp_data[688] = 32'h515fe604;
temp_data[689] = 32'h5160e0c1;
temp_data[690] = 32'h5161d9dc;
temp_data[691] = 32'h5162d196;
temp_data[692] = 32'h5163c836;
temp_data[693] = 32'h5164be16;
temp_data[694] = 32'h5165b392;
temp_data[695] = 32'h5166a911;
temp_data[696] = 32'h51679efe;
temp_data[697] = 32'h516895d1;
temp_data[698] = 32'h51698e0d;
temp_data[699] = 32'h516a883c;
temp_data[700] = 32'h516b84f5;
temp_data[701] = 32'h516c84dc;
temp_data[702] = 32'h516d88a4;
temp_data[703] = 32'h516e9110;
temp_data[704] = 32'h516f9ee9;
temp_data[705] = 32'h5170b31c;
temp_data[706] = 32'h5171ce96;
temp_data[707] = 32'h5172f26f;
temp_data[708] = 32'h51741fcd;
temp_data[709] = 32'h517557f3;
temp_data[710] = 32'h51769c45;
temp_data[711] = 32'h5177ee4a;
temp_data[712] = 32'h51794fb5;
temp_data[713] = 32'h517ac259;
temp_data[714] = 32'h517c4849;
temp_data[715] = 32'h517de3c1;
temp_data[716] = 32'h517f9742;
temp_data[717] = 32'h51816588;
temp_data[718] = 32'h518351a0;
temp_data[719] = 32'h51855eea;
temp_data[720] = 32'h5187911d;
temp_data[721] = 32'h5189ec5f;
temp_data[722] = 32'h518c753a;
temp_data[723] = 32'h518f30c6;
temp_data[724] = 32'h5192249a;
temp_data[725] = 32'h519556eb;
temp_data[726] = 32'h5198ce9e;
temp_data[727] = 32'h519c9353;
temp_data[728] = 32'h51a0ad75;
temp_data[729] = 32'h51a52663;
temp_data[730] = 32'h51aa0870;
temp_data[731] = 32'h51af5f0b;
temp_data[732] = 32'h51b536e3;
temp_data[733] = 32'h51bb9ded;
temp_data[734] = 32'h51c2a3a5;
temp_data[735] = 32'h51ca5921;
temp_data[736] = 32'h51d2d13d;
temp_data[737] = 32'h51dc20cd;
temp_data[738] = 32'h51e65ed5;
temp_data[739] = 32'h51f1a4d3;
temp_data[740] = 32'h51fc37d6;
temp_data[741] = 32'h5205bc7b;
temp_data[742] = 32'h520e4a41;
temp_data[743] = 32'h5215f61f;
temp_data[744] = 32'h521cd2cc;
temp_data[745] = 32'h5222f0d8;
temp_data[746] = 32'h52285ed5;
temp_data[747] = 32'h522d2991;
temp_data[748] = 32'h52315c1c;
temp_data[749] = 32'h5234fff3;
temp_data[750] = 32'h52381d15;
temp_data[751] = 32'h523aba0f;
temp_data[752] = 32'h523cdc1a;
temp_data[753] = 32'h523e871a;
temp_data[754] = 32'h523fbdc2;
temp_data[755] = 32'h52408177;
temp_data[756] = 32'h5240d270;
temp_data[757] = 32'h5240afb8;
temp_data[758] = 32'h52401712;
temp_data[759] = 32'h523f0518;
temp_data[760] = 32'h523d7514;
temp_data[761] = 32'h523b6113;
temp_data[762] = 32'h5238c1b5;
temp_data[763] = 32'h52358e32;
temp_data[764] = 32'h5231bc49;
temp_data[765] = 32'h522d4007;
temp_data[766] = 32'h52280bd4;
temp_data[767] = 32'h5222102c;
temp_data[768] = 32'h521b3b6d;
temp_data[769] = 32'h52154f5d;
temp_data[770] = 32'h52103a79;
temp_data[771] = 32'h520bed74;
temp_data[772] = 32'h52085aee;
temp_data[773] = 32'h5205776c;
temp_data[774] = 32'h52033922;
temp_data[775] = 32'h520197ea;
temp_data[776] = 32'h52008d26;
temp_data[777] = 32'h520013b2;
temp_data[778] = 32'h520027dd;
temp_data[779] = 32'h5200c765;
temp_data[780] = 32'h5201f15a;
temp_data[781] = 32'h5203a63b;
temp_data[782] = 32'h5205e7ef;
temp_data[783] = 32'h5208b9bb;
temp_data[784] = 32'h520c206d;
temp_data[785] = 32'h52102242;
temp_data[786] = 32'h5214c726;
temp_data[787] = 32'h521a18a4;
temp_data[788] = 32'h52202210;
temp_data[789] = 32'h5226f0b7;
temp_data[790] = 32'h522e93e2;
temp_data[791] = 32'h52371d1d;
temp_data[792] = 32'h5240a066;
temp_data[793] = 32'h524b3455;
temp_data[794] = 32'h5256f25a;
temp_data[795] = 32'h5263f71a;
temp_data[796] = 32'h527262a6;
temp_data[797] = 32'h528258d1;
temp_data[798] = 32'h5294019b;
temp_data[799] = 32'h52a78994;
temp_data[800] = 32'h52bd224f;
temp_data[801] = 32'h52d502eb;
temp_data[802] = 32'h52ef688c;
temp_data[803] = 32'h530c970f;
temp_data[804] = 32'h532cd9ae;
temp_data[805] = 32'h535083a9;
temp_data[806] = 32'h5377f139;
temp_data[807] = 32'h53a3885d;
temp_data[808] = 32'h53d3b9e5;
temp_data[809] = 32'h540902c9;
temp_data[810] = 32'h543f598a;
temp_data[811] = 32'h54706d72;
temp_data[812] = 32'h549cbe16;
temp_data[813] = 32'h54c4be83;
temp_data[814] = 32'h54e8d6bb;
temp_data[815] = 32'h550964b6;
temp_data[816] = 32'h5526bd5a;
temp_data[817] = 32'h55412d41;
temp_data[818] = 32'h5558f97f;
temp_data[819] = 32'h556e605f;
temp_data[820] = 32'h558199e1;
temp_data[821] = 32'h5592d86b;
temp_data[822] = 32'h55a24938;
temp_data[823] = 32'h55b014d3;
temp_data[824] = 32'h55bc5f85;
temp_data[825] = 32'h55c749ae;
temp_data[826] = 32'h55d0f01c;
temp_data[827] = 32'h55d96c66;
temp_data[828] = 32'h55e0d524;
temp_data[829] = 32'h55e73e29;
temp_data[830] = 32'h55ecb8d0;
temp_data[831] = 32'h55f15409;
temp_data[832] = 32'h55f51cac;
temp_data[833] = 32'h55f81d75;
temp_data[834] = 32'h55fa5f42;
temp_data[835] = 32'h55fbe914;
temp_data[836] = 32'h55fcc033;
temp_data[837] = 32'h55fce83a;
temp_data[838] = 32'h55fc6313;
temp_data[839] = 32'h55fb3116;
temp_data[840] = 32'h55f950f4;
temp_data[841] = 32'h55f6bfbe;
temp_data[842] = 32'h55f378d9;
temp_data[843] = 32'h55ef75f3;
temp_data[844] = 32'h55eaaef7;
temp_data[845] = 32'h55e519f0;
temp_data[846] = 32'h55deaae3;
temp_data[847] = 32'h55d753c5;
temp_data[848] = 32'h55cf044b;
temp_data[849] = 32'h55c5a9b0;
temp_data[850] = 32'h55bb2e94;
temp_data[851] = 32'h55af7ab7;
temp_data[852] = 32'h55a272b9;
temp_data[853] = 32'h5593f7cf;
temp_data[854] = 32'h5583e775;
temp_data[855] = 32'h55721b09;
temp_data[856] = 32'h555e6773;
temp_data[857] = 32'h55489ca2;
temp_data[858] = 32'h5530851b;
temp_data[859] = 32'h5515e569;
temp_data[860] = 32'h54f87b89;
temp_data[861] = 32'h54d7fe37;
temp_data[862] = 32'h54b41c43;
temp_data[863] = 32'h548c7bc4;
temp_data[864] = 32'h5460b91f;
temp_data[865] = 32'h54306627;
temp_data[866] = 32'h53fb08ff;
temp_data[867] = 32'h53c01a5d;
temp_data[868] = 32'h53888577;
temp_data[869] = 32'h53561d7a;
temp_data[870] = 32'h53286345;
temp_data[871] = 32'h52fee3d6;
temp_data[872] = 32'h52d93726;
temp_data[873] = 32'h52b6ff1e;
temp_data[874] = 32'h5297e697;
temp_data[875] = 32'h527ba09d;
temp_data[876] = 32'h5261e79f;
temp_data[877] = 32'h524a7cbf;
temp_data[878] = 32'h52352735;
temp_data[879] = 32'h5221b3af;
temp_data[880] = 32'h520ff3e9;
temp_data[881] = 32'h51ffbe12;
temp_data[882] = 32'h51f0ec74;
temp_data[883] = 32'h51e35d0b;
temp_data[884] = 32'h51d6f120;
temp_data[885] = 32'h51cb8d09;
temp_data[886] = 32'h51c117c2;
temp_data[887] = 32'h51b77acc;
temp_data[888] = 32'h51aea1d3;
temp_data[889] = 32'h51a67a85;
temp_data[890] = 32'h519ef456;
temp_data[891] = 32'h51980058;
temp_data[892] = 32'h51919121;
temp_data[893] = 32'h518b9a80;
temp_data[894] = 32'h51861188;
temp_data[895] = 32'h5180ec46;
temp_data[896] = 32'h517c21d5;
temp_data[897] = 32'h5177aa19;
temp_data[898] = 32'h51737dcc;
temp_data[899] = 32'h516f964f;
temp_data[900] = 32'h516beda6;
temp_data[901] = 32'h51687e74;
temp_data[902] = 32'h516543d0;
temp_data[903] = 32'h51623950;
temp_data[904] = 32'h515f5aee;
temp_data[905] = 32'h515ca509;
temp_data[906] = 32'h515a1451;
temp_data[907] = 32'h5157a5ca;
temp_data[908] = 32'h515556c1;
temp_data[909] = 32'h515324b7;
temp_data[910] = 32'h51510d6f;
temp_data[911] = 32'h514f0ee0;
temp_data[912] = 32'h514d2731;
temp_data[913] = 32'h514b54a4;
temp_data[914] = 32'h514995bc;
temp_data[915] = 32'h5147e903;
temp_data[916] = 32'h51464d38;
temp_data[917] = 32'h5144c12b;
temp_data[918] = 32'h514343c8;
temp_data[919] = 32'h5141d413;
temp_data[920] = 32'h51407122;
temp_data[921] = 32'h513f1a1e;
temp_data[922] = 32'h513dce4f;
temp_data[923] = 32'h513c8cf4;
temp_data[924] = 32'h513b5571;
temp_data[925] = 32'h513a2728;
temp_data[926] = 32'h51390193;
temp_data[927] = 32'h5137e42a;
temp_data[928] = 32'h5136ce79;
temp_data[929] = 32'h5135c00e;
temp_data[930] = 32'h5134b884;
temp_data[931] = 32'h5133b778;
temp_data[932] = 32'h5132bc99;
temp_data[933] = 32'h5131c78a;
temp_data[934] = 32'h5130d806;
temp_data[935] = 32'h512fedc4;
temp_data[936] = 32'h512f0881;
temp_data[937] = 32'h512e27fa;
temp_data[938] = 32'h512d4bf9;
temp_data[939] = 32'h512c7447;
temp_data[940] = 32'h512ba0ae;
temp_data[941] = 32'h512ad0ff;
temp_data[942] = 32'h512a050c;
temp_data[943] = 32'h51293ca7;
temp_data[944] = 32'h512877af;
temp_data[945] = 32'h5127b5f6;
temp_data[946] = 32'h5126f75e;
temp_data[947] = 32'h51263bc1;
temp_data[948] = 32'h512582fd;
temp_data[949] = 32'h5124ccf7;
temp_data[950] = 32'h5124198f;
temp_data[951] = 32'h512368ad;
temp_data[952] = 32'h5122ba30;
temp_data[953] = 32'h51220e06;
temp_data[954] = 32'h51216413;
temp_data[955] = 32'h5120bc45;
temp_data[956] = 32'h5120167b;
temp_data[957] = 32'h511f72ac;
temp_data[958] = 32'h511ed0bb;
temp_data[959] = 32'h511e309c;
temp_data[960] = 32'h511d923a;
temp_data[961] = 32'h511cf57f;
temp_data[962] = 32'h511c5a64;
temp_data[963] = 32'h511bc0cf;
temp_data[964] = 32'h511b28b3;
temp_data[965] = 32'h511a9204;
temp_data[966] = 32'h5119fcb5;
temp_data[967] = 32'h511968b2;
temp_data[968] = 32'h5118d5f5;
temp_data[969] = 32'h5118446b;
temp_data[970] = 32'h5117b40b;
temp_data[971] = 32'h511724c8;
temp_data[972] = 32'h5116969e;
temp_data[973] = 32'h51160978;
temp_data[974] = 32'h51157d52;
temp_data[975] = 32'h5114f224;
temp_data[976] = 32'h511467e0;
temp_data[977] = 32'h5113de7f;
temp_data[978] = 32'h511355fc;
temp_data[979] = 32'h5112ce4f;
temp_data[980] = 32'h5112476f;
temp_data[981] = 32'h5111c155;
temp_data[982] = 32'h51113c04;
temp_data[983] = 32'h5110b76b;
temp_data[984] = 32'h5110338b;
temp_data[985] = 32'h510fb064;
temp_data[986] = 32'h510f2df1;
temp_data[987] = 32'h510eac32;
temp_data[988] = 32'h510e2b24;
temp_data[989] = 32'h510daac5;
temp_data[990] = 32'h510d2b1b;
temp_data[991] = 32'h510cac26;
temp_data[992] = 32'h510c2de8;
temp_data[993] = 32'h510bb06c;
temp_data[994] = 32'h510b33b9;
temp_data[995] = 32'h510ab7d4;
temp_data[996] = 32'h510a3cc5;
temp_data[997] = 32'h5109c2a0;
temp_data[998] = 32'h51094973;
temp_data[999] = 32'h5108d14a;
temp_data[1000] = 32'h51085a42;
temp_data[1001] = 32'h5107e46d;
temp_data[1002] = 32'h51076fe7;
temp_data[1003] = 32'h5106fcd6;
temp_data[1004] = 32'h51068b54;
temp_data[1005] = 32'h51061b93;
temp_data[1006] = 32'h5105adb8;
temp_data[1007] = 32'h510541ff;
temp_data[1008] = 32'h5104d89d;
temp_data[1009] = 32'h510471da;
temp_data[1010] = 32'h51040dfa;
temp_data[1011] = 32'h5103ad54;
temp_data[1012] = 32'h51035040;
temp_data[1013] = 32'h5102f727;
temp_data[1014] = 32'h5102a283;
temp_data[1015] = 32'h510252d6;
temp_data[1016] = 32'h510208a7;
temp_data[1017] = 32'h5101c4a4;
temp_data[1018] = 32'h5101877b;
temp_data[1019] = 32'h510151f8;
temp_data[1020] = 32'h510124fb;
temp_data[1021] = 32'h51010182;
temp_data[1022] = 32'h5100e8a3;
temp_data[1023] = 32'h5100db90;
temp_data[1024] = 32'h50f714cb;
temp_data[1025] = 32'h50f72114;
temp_data[1026] = 32'h50f7386d;
temp_data[1027] = 32'h50f759a7;
temp_data[1028] = 32'h50f783ae;
temp_data[1029] = 32'h50f7b58d;
temp_data[1030] = 32'h50f7ee63;
temp_data[1031] = 32'h50f82d6b;
temp_data[1032] = 32'h50f871f8;
temp_data[1033] = 32'h50f8bb66;
temp_data[1034] = 32'h50f9092d;
temp_data[1035] = 32'h50f95ac9;
temp_data[1036] = 32'h50f9afc9;
temp_data[1037] = 32'h50fa07c8;
temp_data[1038] = 32'h50fa626b;
temp_data[1039] = 32'h50fabf5d;
temp_data[1040] = 32'h50fb1e5c;
temp_data[1041] = 32'h50fb7f24;
temp_data[1042] = 32'h50fbe17a;
temp_data[1043] = 32'h50fc452c;
temp_data[1044] = 32'h50fcaa0d;
temp_data[1045] = 32'h50fd0ff1;
temp_data[1046] = 32'h50fd76b8;
temp_data[1047] = 32'h50fdde3c;
temp_data[1048] = 32'h50fe4667;
temp_data[1049] = 32'h50feaf21;
temp_data[1050] = 32'h50ff1850;
temp_data[1051] = 32'h50ff81e0;
temp_data[1052] = 32'h50ffebc0;
temp_data[1053] = 32'h510055e7;
temp_data[1054] = 32'h5100c044;
temp_data[1055] = 32'h51012acc;
temp_data[1056] = 32'h51019579;
temp_data[1057] = 32'h5102003b;
temp_data[1058] = 32'h51026b16;
temp_data[1059] = 32'h5102d5fe;
temp_data[1060] = 32'h510340ee;
temp_data[1061] = 32'h5103abe2;
temp_data[1062] = 32'h510416df;
temp_data[1063] = 32'h510481d8;
temp_data[1064] = 32'h5104ecd5;
temp_data[1065] = 32'h510557cd;
temp_data[1066] = 32'h5105c2c6;
temp_data[1067] = 32'h51062dba;
temp_data[1068] = 32'h510698b3;
temp_data[1069] = 32'h510703a7;
temp_data[1070] = 32'h51076ea0;
temp_data[1071] = 32'h5107d99d;
temp_data[1072] = 32'h5108449e;
temp_data[1073] = 32'h5108afa7;
temp_data[1074] = 32'h51091ab9;
temp_data[1075] = 32'h510985d7;
temp_data[1076] = 32'h5109f106;
temp_data[1077] = 32'h510a5c46;
temp_data[1078] = 32'h510ac79b;
temp_data[1079] = 32'h510b330d;
temp_data[1080] = 32'h510b9e95;
temp_data[1081] = 32'h510c0a42;
temp_data[1082] = 32'h510c7610;
temp_data[1083] = 32'h510ce204;
temp_data[1084] = 32'h510d4e23;
temp_data[1085] = 32'h510dba6f;
temp_data[1086] = 32'h510e26f2;
temp_data[1087] = 32'h510e93a7;
temp_data[1088] = 32'h510f009b;
temp_data[1089] = 32'h510f6dca;
temp_data[1090] = 32'h510fdb40;
temp_data[1091] = 32'h511048fe;
temp_data[1092] = 32'h5110b702;
temp_data[1093] = 32'h5111255f;
temp_data[1094] = 32'h5111940c;
temp_data[1095] = 32'h51120315;
temp_data[1096] = 32'h5112727e;
temp_data[1097] = 32'h5112e24c;
temp_data[1098] = 32'h51135283;
temp_data[1099] = 32'h5113c322;
temp_data[1100] = 32'h5114343b;
temp_data[1101] = 32'h5114a5ca;
temp_data[1102] = 32'h511517d7;
temp_data[1103] = 32'h51158a65;
temp_data[1104] = 32'h5115fd7e;
temp_data[1105] = 32'h51167126;
temp_data[1106] = 32'h5116e560;
temp_data[1107] = 32'h51175a36;
temp_data[1108] = 32'h5117cfab;
temp_data[1109] = 32'h511845c8;
temp_data[1110] = 32'h5118bc94;
temp_data[1111] = 32'h51193411;
temp_data[1112] = 32'h5119ac4b;
temp_data[1113] = 32'h511a2546;
temp_data[1114] = 32'h511a9f0a;
temp_data[1115] = 32'h511b19a0;
temp_data[1116] = 32'h511b9510;
temp_data[1117] = 32'h511c115e;
temp_data[1118] = 32'h511c8e93;
temp_data[1119] = 32'h511d0cbb;
temp_data[1120] = 32'h511d8bdf;
temp_data[1121] = 32'h511e0c02;
temp_data[1122] = 32'h511e8d37;
temp_data[1123] = 32'h511f0f80;
temp_data[1124] = 32'h511f92ea;
temp_data[1125] = 32'h51201783;
temp_data[1126] = 32'h51209d52;
temp_data[1127] = 32'h51212464;
temp_data[1128] = 32'h5121acc5;
temp_data[1129] = 32'h51223682;
temp_data[1130] = 32'h5122c1a9;
temp_data[1131] = 32'h51234e44;
temp_data[1132] = 32'h5123dc6a;
temp_data[1133] = 32'h51246c22;
temp_data[1134] = 32'h5124fd82;
temp_data[1135] = 32'h51259097;
temp_data[1136] = 32'h51262574;
temp_data[1137] = 32'h5126bc2c;
temp_data[1138] = 32'h512754d2;
temp_data[1139] = 32'h5127ef78;
temp_data[1140] = 32'h51288c37;
temp_data[1141] = 32'h51292b1f;
temp_data[1142] = 32'h5129cc4b;
temp_data[1143] = 32'h512a6fd6;
temp_data[1144] = 32'h512b15d3;
temp_data[1145] = 32'h512bbe59;
temp_data[1146] = 32'h512c698c;
temp_data[1147] = 32'h512d1783;
temp_data[1148] = 32'h512dc85c;
temp_data[1149] = 32'h512e7c31;
temp_data[1150] = 32'h512f331e;
temp_data[1151] = 32'h512fed4a;
temp_data[1152] = 32'h5130aace;
temp_data[1153] = 32'h51316bc6;
temp_data[1154] = 32'h51323055;
temp_data[1155] = 32'h5132f894;
temp_data[1156] = 32'h5133c4a8;
temp_data[1157] = 32'h513494ab;
temp_data[1158] = 32'h513568b2;
temp_data[1159] = 32'h513640dd;
temp_data[1160] = 32'h51371d3b;
temp_data[1161] = 32'h5137fddf;
temp_data[1162] = 32'h5138e2d6;
temp_data[1163] = 32'h5139cc25;
temp_data[1164] = 32'h513ab9d4;
temp_data[1165] = 32'h513babd6;
temp_data[1166] = 32'h513ca21f;
temp_data[1167] = 32'h513d9c91;
temp_data[1168] = 32'h513e9b0b;
temp_data[1169] = 32'h513f9d5e;
temp_data[1170] = 32'h5140a348;
temp_data[1171] = 32'h5141ac7e;
temp_data[1172] = 32'h5142b89d;
temp_data[1173] = 32'h5143c73f;
temp_data[1174] = 32'h5144d7e4;
temp_data[1175] = 32'h5145e9f7;
temp_data[1176] = 32'h5146fcdb;
temp_data[1177] = 32'h51480fdc;
temp_data[1178] = 32'h5149223a;
temp_data[1179] = 32'h514a3322;
temp_data[1180] = 32'h514b41bc;
temp_data[1181] = 32'h514c4ead;
temp_data[1182] = 32'h514d5f89;
temp_data[1183] = 32'h514e7360;
temp_data[1184] = 32'h514f8961;
temp_data[1185] = 32'h5150a0c7;
temp_data[1186] = 32'h5151b8d8;
temp_data[1187] = 32'h5152d0f2;
temp_data[1188] = 32'h5153e881;
temp_data[1189] = 32'h5154ff09;
temp_data[1190] = 32'h5156141f;
temp_data[1191] = 32'h51572763;
temp_data[1192] = 32'h51583897;
temp_data[1193] = 32'h5159477c;
temp_data[1194] = 32'h515a53f4;
temp_data[1195] = 32'h515b5dea;
temp_data[1196] = 32'h515c654d;
temp_data[1197] = 32'h515d6a2f;
temp_data[1198] = 32'h515e6c9c;
temp_data[1199] = 32'h515f6cb1;
temp_data[1200] = 32'h51606a9c;
temp_data[1201] = 32'h5161668c;
temp_data[1202] = 32'h516260bb;
temp_data[1203] = 32'h51635975;
temp_data[1204] = 32'h51645101;
temp_data[1205] = 32'h516547b6;
temp_data[1206] = 32'h51663df7;
temp_data[1207] = 32'h51673422;
temp_data[1208] = 32'h51682ab2;
temp_data[1209] = 32'h51692214;
temp_data[1210] = 32'h516a1ad6;
temp_data[1211] = 32'h516b157b;
temp_data[1212] = 32'h516c129d;
temp_data[1213] = 32'h516d12e0;
temp_data[1214] = 32'h516e16f8;
temp_data[1215] = 32'h516f1fa7;
temp_data[1216] = 32'h51702dba;
temp_data[1217] = 32'h51714214;
temp_data[1218] = 32'h51725db3;
temp_data[1219] = 32'h5173819d;
temp_data[1220] = 32'h5174aeff;
temp_data[1221] = 32'h5175e721;
temp_data[1222] = 32'h51772b5e;
temp_data[1223] = 32'h51787d41;
temp_data[1224] = 32'h5179de76;
temp_data[1225] = 32'h517b50db;
temp_data[1226] = 32'h517cd673;
temp_data[1227] = 32'h517e7186;
temp_data[1228] = 32'h51802489;
temp_data[1229] = 32'h5181f241;
temp_data[1230] = 32'h5183ddb1;
temp_data[1231] = 32'h5185ea3a;
temp_data[1232] = 32'h51881b8f;
temp_data[1233] = 32'h518a75da;
temp_data[1234] = 32'h518cfda0;
temp_data[1235] = 32'h518fb7f1;
temp_data[1236] = 32'h5192aa6d;
temp_data[1237] = 32'h5195db40;
temp_data[1238] = 32'h51995155;
temp_data[1239] = 32'h519d1440;
temp_data[1240] = 32'h51a12c73;
temp_data[1241] = 32'h51a5a34d;
temp_data[1242] = 32'h51aa831b;
temp_data[1243] = 32'h51afd75a;
temp_data[1244] = 32'h51b5acac;
temp_data[1245] = 32'h51bc1112;
temp_data[1246] = 32'h51c3140a;
temp_data[1247] = 32'h51cac6b0;
temp_data[1248] = 32'h51d33be2;
temp_data[1249] = 32'h51dc887f;
temp_data[1250] = 32'h51e6c38b;
temp_data[1251] = 32'h51f20692;
temp_data[1252] = 32'h51fc96ab;
temp_data[1253] = 32'h52061876;
temp_data[1254] = 32'h520ea37b;
temp_data[1255] = 32'h52164cbe;
temp_data[1256] = 32'h521d26f2;
temp_data[1257] = 32'h522342af;
temp_data[1258] = 32'h5228ae8e;
temp_data[1259] = 32'h522d775c;
temp_data[1260] = 32'h5231a82f;
temp_data[1261] = 32'h52354a84;
temp_data[1262] = 32'h5238665a;
temp_data[1263] = 32'h523b023a;
temp_data[1264] = 32'h523d2360;
temp_data[1265] = 32'h523ecdb3;
temp_data[1266] = 32'h524003da;
temp_data[1267] = 32'h5240c73b;
temp_data[1268] = 32'h5241180d;
temp_data[1269] = 32'h5240f556;
temp_data[1270] = 32'h52405cd5;
temp_data[1271] = 32'h523f4b23;
temp_data[1272] = 32'h523dbb88;
temp_data[1273] = 32'h523ba805;
temp_data[1274] = 32'h5239093e;
temp_data[1275] = 32'h5235d667;
temp_data[1276] = 32'h5232053a;
temp_data[1277] = 32'h522d89c2;
temp_data[1278] = 32'h52285660;
temp_data[1279] = 32'h52225b8a;
temp_data[1280] = 32'h521b87a5;
temp_data[1281] = 32'h52159c6b;
temp_data[1282] = 32'h52108855;
temp_data[1283] = 32'h520c3c10;
temp_data[1284] = 32'h5208aa43;
temp_data[1285] = 32'h5205c765;
temp_data[1286] = 32'h520389ad;
temp_data[1287] = 32'h5201e8e6;
temp_data[1288] = 32'h5200de76;
temp_data[1289] = 32'h52006534;
temp_data[1290] = 32'h5200796c;
temp_data[1291] = 32'h520118ce;
temp_data[1292] = 32'h52024274;
temp_data[1293] = 32'h5203f6cb;
temp_data[1294] = 32'h520637b9;
temp_data[1295] = 32'h52090881;
temp_data[1296] = 32'h520c6ddf;
temp_data[1297] = 32'h52106e1a;
temp_data[1298] = 32'h52151106;
temp_data[1299] = 32'h521a6031;
temp_data[1300] = 32'h522066ed;
temp_data[1301] = 32'h5227326e;
temp_data[1302] = 32'h522ed203;
temp_data[1303] = 32'h5237572a;
temp_data[1304] = 32'h5240d5d8;
temp_data[1305] = 32'h524b649d;
temp_data[1306] = 32'h52571ce3;
temp_data[1307] = 32'h52641b48;
temp_data[1308] = 32'h52727fcc;
temp_data[1309] = 32'h52826e44;
temp_data[1310] = 32'h52940eaa;
temp_data[1311] = 32'h52a78d8f;
temp_data[1312] = 32'h52bd1c82;
temp_data[1313] = 32'h52d4f29d;
temp_data[1314] = 32'h52ef4d16;
temp_data[1315] = 32'h530c6fd2;
temp_data[1316] = 32'h532ca609;
temp_data[1317] = 32'h5350431c;
temp_data[1318] = 32'h5377a351;
temp_data[1319] = 32'h53a32cc3;
temp_data[1320] = 32'h53d35050;
temp_data[1321] = 32'h54088b1a;
temp_data[1322] = 32'h543ed3b3;
temp_data[1323] = 32'h546fd98c;
temp_data[1324] = 32'h549c1c54;
temp_data[1325] = 32'h54c40f34;
temp_data[1326] = 32'h54e81a3f;
temp_data[1327] = 32'h55089b89;
temp_data[1328] = 32'h5525e804;
temp_data[1329] = 32'h55404c59;
temp_data[1330] = 32'h55580dae;
temp_data[1331] = 32'h556d6a44;
temp_data[1332] = 32'h55809a31;
temp_data[1333] = 32'h5591cfcc;
temp_data[1334] = 32'h55a13854;
temp_data[1335] = 32'h55aefc54;
temp_data[1336] = 32'h55bb4007;
temp_data[1337] = 32'h55c623c8;
temp_data[1338] = 32'h55cfc469;
temp_data[1339] = 32'h55d83b71;
temp_data[1340] = 32'h55df9f6f;
temp_data[1341] = 32'h55e60432;
temp_data[1342] = 32'h55eb7b0b;
temp_data[1343] = 32'h55f012e8;
temp_data[1344] = 32'h55f3d895;
temp_data[1345] = 32'h55f6d6d0;
temp_data[1346] = 32'h55f9166e;
temp_data[1347] = 32'h55fa9e6b;
temp_data[1348] = 32'h55fb7410;
temp_data[1349] = 32'h55fb9af2;
temp_data[1350] = 32'h55fb14fd;
temp_data[1351] = 32'h55f9e282;
temp_data[1352] = 32'h55f8023a;
temp_data[1353] = 32'h55f57132;
temp_data[1354] = 32'h55f22ad4;
temp_data[1355] = 32'h55ee28d0;
temp_data[1356] = 32'h55e9630f;
temp_data[1357] = 32'h55e3cfa7;
temp_data[1358] = 32'h55dd629e;
temp_data[1359] = 32'h55d60df6;
temp_data[1360] = 32'h55cdc161;
temp_data[1361] = 32'h55c46a2b;
temp_data[1362] = 32'h55b9f2f1;
temp_data[1363] = 32'h55ae437c;
temp_data[1364] = 32'h55a14079;
temp_data[1365] = 32'h5592cb21;
temp_data[1366] = 32'h5582c0f4;
temp_data[1367] = 32'h5570fb5d;
temp_data[1368] = 32'h555d4f3c;
temp_data[1369] = 32'h55478c8b;
temp_data[1370] = 32'h552f7dcc;
temp_data[1371] = 32'h5514e786;
temp_data[1372] = 32'h54f787b1;
temp_data[1373] = 32'h54d71501;
temp_data[1374] = 32'h54b33e36;
temp_data[1375] = 32'h548ba954;
temp_data[1376] = 32'h545ff2b2;
temp_data[1377] = 32'h542fac08;
temp_data[1378] = 32'h53fa5b5b;
temp_data[1379] = 32'h53bf794a;
temp_data[1380] = 32'h5387f0ed;
temp_data[1381] = 32'h5355955b;
temp_data[1382] = 32'h5327e74f;
temp_data[1383] = 32'h52fe73b4;
temp_data[1384] = 32'h52d8d274;
temp_data[1385] = 32'h52b6a555;
temp_data[1386] = 32'h52979731;
temp_data[1387] = 32'h527b5b08;
temp_data[1388] = 32'h5261ab36;
temp_data[1389] = 32'h524a48e4;
temp_data[1390] = 32'h5234fb40;
temp_data[1391] = 32'h52218f04;
temp_data[1392] = 32'h520fd5e9;
temp_data[1393] = 32'h51ffa62b;
temp_data[1394] = 32'h51f0da12;
temp_data[1395] = 32'h51e34fa9;
temp_data[1396] = 32'h51d6e83e;
temp_data[1397] = 32'h51cb882b;
temp_data[1398] = 32'h51c11683;
temp_data[1399] = 32'h51b77cbf;
temp_data[1400] = 32'h51aea6a0;
temp_data[1401] = 32'h51a681d4;
temp_data[1402] = 32'h519efddb;
temp_data[1403] = 32'h51980bd0;
temp_data[1404] = 32'h51919e49;
temp_data[1405] = 32'h518ba922;
temp_data[1406] = 32'h5186216c;
temp_data[1407] = 32'h5180fd48;
temp_data[1408] = 32'h517c33c2;
temp_data[1409] = 32'h5177bcd3;
temp_data[1410] = 32'h5173912e;
temp_data[1411] = 32'h516faa3b;
temp_data[1412] = 32'h516c0208;
temp_data[1413] = 32'h51689332;
temp_data[1414] = 32'h516558d6;
temp_data[1415] = 32'h51624e8b;
temp_data[1416] = 32'h515f704c;
temp_data[1417] = 32'h515cba7c;
temp_data[1418] = 32'h515a29d0;
temp_data[1419] = 32'h5157bb49;
temp_data[1420] = 32'h51556c33;
temp_data[1421] = 32'h51533a19;
temp_data[1422] = 32'h515122b8;
temp_data[1423] = 32'h514f2407;
temp_data[1424] = 32'h514d3c2e;
temp_data[1425] = 32'h514b697b;
temp_data[1426] = 32'h5149aa61;
temp_data[1427] = 32'h5147fd76;
temp_data[1428] = 32'h51466174;
temp_data[1429] = 32'h5144d530;
temp_data[1430] = 32'h5143578e;
temp_data[1431] = 32'h5141e79b;
temp_data[1432] = 32'h5140846a;
temp_data[1433] = 32'h513f2d2c;
temp_data[1434] = 32'h513de115;
temp_data[1435] = 32'h513c9f7b;
temp_data[1436] = 32'h513b67b2;
temp_data[1437] = 32'h513a392a;
temp_data[1438] = 32'h5139134d;
temp_data[1439] = 32'h5137f5a1;
temp_data[1440] = 32'h5136dfa8;
temp_data[1441] = 32'h5135d0fa;
temp_data[1442] = 32'h5134c92a;
temp_data[1443] = 32'h5133c7de;
temp_data[1444] = 32'h5132ccb8;
temp_data[1445] = 32'h5131d767;
temp_data[1446] = 32'h5130e79f;
temp_data[1447] = 32'h512ffd1a;
temp_data[1448] = 32'h512f178f;
temp_data[1449] = 32'h512e36ca;
temp_data[1450] = 32'h512d5a86;
temp_data[1451] = 32'h512c8290;
temp_data[1452] = 32'h512baeb4;
temp_data[1453] = 32'h512adec6;
temp_data[1454] = 32'h512a1290;
temp_data[1455] = 32'h512949ed;
temp_data[1456] = 32'h512884b6;
temp_data[1457] = 32'h5127c2bd;
temp_data[1458] = 32'h512703e6;
temp_data[1459] = 32'h5126480a;
temp_data[1460] = 32'h51258f08;
temp_data[1461] = 32'h5124d8c7;
temp_data[1462] = 32'h51242520;
temp_data[1463] = 32'h51237400;
temp_data[1464] = 32'h5122c54c;
temp_data[1465] = 32'h512218e7;
temp_data[1466] = 32'h51216eb9;
temp_data[1467] = 32'h5120c6ac;
temp_data[1468] = 32'h512020ab;
temp_data[1469] = 32'h511f7ca2;
temp_data[1470] = 32'h511eda77;
temp_data[1471] = 32'h511e3a21;
temp_data[1472] = 32'h511d9b84;
temp_data[1473] = 32'h511cfe93;
temp_data[1474] = 32'h511c633d;
temp_data[1475] = 32'h511bc971;
temp_data[1476] = 32'h511b3123;
temp_data[1477] = 32'h511a9a3d;
temp_data[1478] = 32'h511a04b8;
temp_data[1479] = 32'h5119707e;
temp_data[1480] = 32'h5118dd8b;
temp_data[1481] = 32'h51184bcf;
temp_data[1482] = 32'h5117bb38;
temp_data[1483] = 32'h51172bc3;
temp_data[1484] = 32'h51169d62;
temp_data[1485] = 32'h5116100a;
temp_data[1486] = 32'h511583b2;
temp_data[1487] = 32'h5114f851;
temp_data[1488] = 32'h51146ddb;
temp_data[1489] = 32'h5113e447;
temp_data[1490] = 32'h51135b92;
temp_data[1491] = 32'h5112d3b3;
temp_data[1492] = 32'h51124ca5;
temp_data[1493] = 32'h5111c65c;
temp_data[1494] = 32'h511140d5;
temp_data[1495] = 32'h5110bc0e;
temp_data[1496] = 32'h51103800;
temp_data[1497] = 32'h510fb4ab;
temp_data[1498] = 32'h510f3209;
temp_data[1499] = 32'h510eb018;
temp_data[1500] = 32'h510e2ed8;
temp_data[1501] = 32'h510dae4b;
temp_data[1502] = 32'h510d2e73;
temp_data[1503] = 32'h510caf53;
temp_data[1504] = 32'h510c30e8;
temp_data[1505] = 32'h510bb342;
temp_data[1506] = 32'h510b3661;
temp_data[1507] = 32'h510aba4d;
temp_data[1508] = 32'h510a3f14;
temp_data[1509] = 32'h5109c4c6;
temp_data[1510] = 32'h51094b6a;
temp_data[1511] = 32'h5108d317;
temp_data[1512] = 32'h51085be6;
temp_data[1513] = 32'h5107e5e6;
temp_data[1514] = 32'h5107713b;
temp_data[1515] = 32'h5106fdfc;
temp_data[1516] = 32'h51068c54;
temp_data[1517] = 32'h51061c6d;
temp_data[1518] = 32'h5105ae6d;
temp_data[1519] = 32'h5105428d;
temp_data[1520] = 32'h5104d90a;
temp_data[1521] = 32'h51047222;
temp_data[1522] = 32'h51040e1b;
temp_data[1523] = 32'h5103ad54;
temp_data[1524] = 32'h5103501e;
temp_data[1525] = 32'h5102f6ec;
temp_data[1526] = 32'h5102a227;
temp_data[1527] = 32'h5102525d;
temp_data[1528] = 32'h51020818;
temp_data[1529] = 32'h5101c3f8;
temp_data[1530] = 32'h510186ba;
temp_data[1531] = 32'h51015126;
temp_data[1532] = 32'h51012418;
temp_data[1533] = 32'h51010093;
temp_data[1534] = 32'h5100e7a7;
temp_data[1535] = 32'h5100da94;
temp_data[1536] = 32'h50f70e6f;
temp_data[1537] = 32'h50f71abd;
temp_data[1538] = 32'h50f7321e;
temp_data[1539] = 32'h50f75369;
temp_data[1540] = 32'h50f77d80;
temp_data[1541] = 32'h50f7af71;
temp_data[1542] = 32'h50f7e860;
temp_data[1543] = 32'h50f82785;
temp_data[1544] = 32'h50f86c2f;
temp_data[1545] = 32'h50f8b5bf;
temp_data[1546] = 32'h50f903a3;
temp_data[1547] = 32'h50f95565;
temp_data[1548] = 32'h50f9aa8b;
temp_data[1549] = 32'h50fa02b0;
temp_data[1550] = 32'h50fa5d7d;
temp_data[1551] = 32'h50faba9d;
temp_data[1552] = 32'h50fb19c6;
temp_data[1553] = 32'h50fb7abc;
temp_data[1554] = 32'h50fbdd40;
temp_data[1555] = 32'h50fc4120;
temp_data[1556] = 32'h50fca62f;
temp_data[1557] = 32'h50fd0c46;
temp_data[1558] = 32'h50fd733b;
temp_data[1559] = 32'h50fddaf5;
temp_data[1560] = 32'h50fe4352;
temp_data[1561] = 32'h50feac3f;
temp_data[1562] = 32'h50ff15a0;
temp_data[1563] = 32'h50ff7f63;
temp_data[1564] = 32'h50ffe97d;
temp_data[1565] = 32'h510053d6;
temp_data[1566] = 32'h5100be6a;
temp_data[1567] = 32'h51012928;
temp_data[1568] = 32'h51019408;
temp_data[1569] = 32'h5101ff04;
temp_data[1570] = 32'h51026a12;
temp_data[1571] = 32'h5102d530;
temp_data[1572] = 32'h5103405b;
temp_data[1573] = 32'h5103ab8a;
temp_data[1574] = 32'h510416b9;
temp_data[1575] = 32'h510481ed;
temp_data[1576] = 32'h5104ed20;
temp_data[1577] = 32'h51055853;
temp_data[1578] = 32'h5105c387;
temp_data[1579] = 32'h51062eb6;
temp_data[1580] = 32'h510699e5;
temp_data[1581] = 32'h51070514;
temp_data[1582] = 32'h51077048;
temp_data[1583] = 32'h5107db7f;
temp_data[1584] = 32'h510846bb;
temp_data[1585] = 32'h5108b1ff;
temp_data[1586] = 32'h51091d4b;
temp_data[1587] = 32'h510988a4;
temp_data[1588] = 32'h5109f40e;
temp_data[1589] = 32'h510a5f8d;
temp_data[1590] = 32'h510acb1d;
temp_data[1591] = 32'h510b36ca;
temp_data[1592] = 32'h510ba290;
temp_data[1593] = 32'h510c0e78;
temp_data[1594] = 32'h510c7a85;
temp_data[1595] = 32'h510ce6b4;
temp_data[1596] = 32'h510d5311;
temp_data[1597] = 32'h510dbf9c;
temp_data[1598] = 32'h510e2c5e;
temp_data[1599] = 32'h510e9952;
temp_data[1600] = 32'h510f0685;
temp_data[1601] = 32'h510f73f3;
temp_data[1602] = 32'h510fe1a8;
temp_data[1603] = 32'h51104fa5;
temp_data[1604] = 32'h5110bdec;
temp_data[1605] = 32'h51112c88;
temp_data[1606] = 32'h51119b78;
temp_data[1607] = 32'h51120ac4;
temp_data[1608] = 32'h51127a70;
temp_data[1609] = 32'h5112ea7d;
temp_data[1610] = 32'h51135af7;
temp_data[1611] = 32'h5113cbda;
temp_data[1612] = 32'h51143d36;
temp_data[1613] = 32'h5114af08;
temp_data[1614] = 32'h51152157;
temp_data[1615] = 32'h5115942d;
temp_data[1616] = 32'h5116078e;
temp_data[1617] = 32'h51167b78;
temp_data[1618] = 32'h5116effe;
temp_data[1619] = 32'h5117651b;
temp_data[1620] = 32'h5117dad7;
temp_data[1621] = 32'h51185140;
temp_data[1622] = 32'h5118c854;
temp_data[1623] = 32'h5119401c;
temp_data[1624] = 32'h5119b8a2;
temp_data[1625] = 32'h511a31e8;
temp_data[1626] = 32'h511aabfc;
temp_data[1627] = 32'h511b26dd;
temp_data[1628] = 32'h511ba298;
temp_data[1629] = 32'h511c1f36;
temp_data[1630] = 32'h511c9cbf;
temp_data[1631] = 32'h511d1b3b;
temp_data[1632] = 32'h511d9aae;
temp_data[1633] = 32'h511e1b2a;
temp_data[1634] = 32'h511e9cb2;
temp_data[1635] = 32'h511f1f4f;
temp_data[1636] = 32'h511fa316;
temp_data[1637] = 32'h51202807;
temp_data[1638] = 32'h5120ae2e;
temp_data[1639] = 32'h512135a0;
temp_data[1640] = 32'h5121be5e;
temp_data[1641] = 32'h5122487c;
temp_data[1642] = 32'h5122d406;
temp_data[1643] = 32'h5123610b;
temp_data[1644] = 32'h5123ef95;
temp_data[1645] = 32'h51247fbb;
temp_data[1646] = 32'h51251188;
temp_data[1647] = 32'h5125a512;
temp_data[1648] = 32'h51263a64;
temp_data[1649] = 32'h5126d191;
temp_data[1650] = 32'h51276ab6;
temp_data[1651] = 32'h512805de;
temp_data[1652] = 32'h5128a323;
temp_data[1653] = 32'h51294296;
temp_data[1654] = 32'h5129e454;
temp_data[1655] = 32'h512a8876;
temp_data[1656] = 32'h512b2f12;
temp_data[1657] = 32'h512bd845;
temp_data[1658] = 32'h512c8427;
temp_data[1659] = 32'h512d32d7;
temp_data[1660] = 32'h512de475;
temp_data[1661] = 32'h512e991c;
temp_data[1662] = 32'h512f50e7;
temp_data[1663] = 32'h51300bfe;
temp_data[1664] = 32'h5130ca7d;
temp_data[1665] = 32'h51318c82;
temp_data[1666] = 32'h51325233;
temp_data[1667] = 32'h51331bac;
temp_data[1668] = 32'h5133e90c;
temp_data[1669] = 32'h5134ba73;
temp_data[1670] = 32'h51359000;
temp_data[1671] = 32'h513669cb;
temp_data[1672] = 32'h513747ed;
temp_data[1673] = 32'h51382a7c;
temp_data[1674] = 32'h51391184;
temp_data[1675] = 32'h5139fd11;
temp_data[1676] = 32'h513aed29;
temp_data[1677] = 32'h513be1ca;
temp_data[1678] = 32'h513cdae4;
temp_data[1679] = 32'h513dd862;
temp_data[1680] = 32'h513eda23;
temp_data[1681] = 32'h513fdff4;
temp_data[1682] = 32'h5140e99f;
temp_data[1683] = 32'h5141f6d3;
temp_data[1684] = 32'h51430731;
temp_data[1685] = 32'h51441a4c;
temp_data[1686] = 32'h51452fa5;
temp_data[1687] = 32'h514646a6;
temp_data[1688] = 32'h51475ea6;
temp_data[1689] = 32'h514876ee;
temp_data[1690] = 32'h51498eb4;
temp_data[1691] = 32'h514aa51e;
temp_data[1692] = 32'h514bb941;
temp_data[1693] = 32'h514ccbc9;
temp_data[1694] = 32'h514de22a;
temp_data[1695] = 32'h514efb7a;
temp_data[1696] = 32'h515016d3;
temp_data[1697] = 32'h5151336e;
temp_data[1698] = 32'h51525083;
temp_data[1699] = 32'h51536d6e;
temp_data[1700] = 32'h51548998;
temp_data[1701] = 32'h5155a47b;
temp_data[1702] = 32'h5156bdad;
temp_data[1703] = 32'h5157d4d0;
temp_data[1704] = 32'h5158e99f;
temp_data[1705] = 32'h5159fbe7;
temp_data[1706] = 32'h515b0b80;
temp_data[1707] = 32'h515c1859;
temp_data[1708] = 32'h515d226c;
temp_data[1709] = 32'h515e29c7;
temp_data[1710] = 32'h515f2e77;
temp_data[1711] = 32'h516030a5;
temp_data[1712] = 32'h5161307b;
temp_data[1713] = 32'h51622e2c;
temp_data[1714] = 32'h516329fa;
temp_data[1715] = 32'h5164242d;
temp_data[1716] = 32'h51651d11;
temp_data[1717] = 32'h51661501;
temp_data[1718] = 32'h51670c5f;
temp_data[1719] = 32'h51680392;
temp_data[1720] = 32'h5168fb0d;
temp_data[1721] = 32'h5169f345;
temp_data[1722] = 32'h516aecc4;
temp_data[1723] = 32'h516be810;
temp_data[1724] = 32'h516ce5cd;
temp_data[1725] = 32'h516de697;
temp_data[1726] = 32'h516eeb20;
temp_data[1727] = 32'h516ff42c;
temp_data[1728] = 32'h5171028e;
temp_data[1729] = 32'h51721722;
temp_data[1730] = 32'h517332ec;
temp_data[1731] = 32'h517456ef;
temp_data[1732] = 32'h51758455;
temp_data[1733] = 32'h5176bc62;
temp_data[1734] = 32'h5178007a;
temp_data[1735] = 32'h51795226;
temp_data[1736] = 32'h517ab307;
temp_data[1737] = 32'h517c2503;
temp_data[1738] = 32'h517daa19;
temp_data[1739] = 32'h517f4489;
temp_data[1740] = 32'h5180f6cb;
temp_data[1741] = 32'h5182c3a0;
temp_data[1742] = 32'h5184ae10;
temp_data[1743] = 32'h5186b96f;
temp_data[1744] = 32'h5188e975;
temp_data[1745] = 32'h518b4242;
temp_data[1746] = 32'h518dc85c;
temp_data[1747] = 32'h519080d4;
temp_data[1748] = 32'h5193713f;
temp_data[1749] = 32'h51969fcf;
temp_data[1750] = 32'h519a1362;
temp_data[1751] = 32'h519dd399;
temp_data[1752] = 32'h51a1e8d9;
temp_data[1753] = 32'h51a65c85;
temp_data[1754] = 32'h51ab38eb;
temp_data[1755] = 32'h51b08983;
temp_data[1756] = 32'h51b65afb;
temp_data[1757] = 32'h51bcbb5a;
temp_data[1758] = 32'h51c3ba1b;
temp_data[1759] = 32'h51cb6862;
temp_data[1760] = 32'h51d3d91f;
temp_data[1761] = 32'h51dd2132;
temp_data[1762] = 32'h51e757b0;
temp_data[1763] = 32'h51f29629;
temp_data[1764] = 32'h51fd21c9;
temp_data[1765] = 32'h52069f34;
temp_data[1766] = 32'h520f2603;
temp_data[1767] = 32'h5216cb3e;
temp_data[1768] = 32'h521da1a5;
temp_data[1769] = 32'h5223b9d8;
temp_data[1770] = 32'h52292279;
temp_data[1771] = 32'h522de853;
temp_data[1772] = 32'h52321683;
temp_data[1773] = 32'h5235b689;
temp_data[1774] = 32'h5238d05f;
temp_data[1775] = 32'h523b6a94;
temp_data[1776] = 32'h523d8a59;
temp_data[1777] = 32'h523f339c;
temp_data[1778] = 32'h524068f9;
temp_data[1779] = 32'h52412bdc;
temp_data[1780] = 32'h52417c70;
temp_data[1781] = 32'h524159b4;
temp_data[1782] = 32'h5240c16a;
temp_data[1783] = 32'h523fb021;
temp_data[1784] = 32'h523e211d;
temp_data[1785] = 32'h523c0e5a;
temp_data[1786] = 32'h5239707a;
temp_data[1787] = 32'h52363ea3;
temp_data[1788] = 32'h52326e8f;
temp_data[1789] = 32'h522df445;
temp_data[1790] = 32'h5228c21a;
temp_data[1791] = 32'h5222c886;
temp_data[1792] = 32'h521bf5e0;
temp_data[1793] = 32'h52160be5;
temp_data[1794] = 32'h5210f909;
temp_data[1795] = 32'h520cadeb;
temp_data[1796] = 32'h52091d2e;
temp_data[1797] = 32'h52063b47;
temp_data[1798] = 32'h5203fe61;
temp_data[1799] = 32'h52025e46;
temp_data[1800] = 32'h52015454;
temp_data[1801] = 32'h5200db5e;
temp_data[1802] = 32'h5200efa2;
temp_data[1803] = 32'h52018ece;
temp_data[1804] = 32'h5202b7f1;
temp_data[1805] = 32'h52046b76;
temp_data[1806] = 32'h5206ab36;
temp_data[1807] = 32'h52097a6c;
temp_data[1808] = 32'h520cddce;
temp_data[1809] = 32'h5210db90;
temp_data[1810] = 32'h52157b89;
temp_data[1811] = 32'h521ac732;
temp_data[1812] = 32'h5220c9d1;
temp_data[1813] = 32'h52279093;
temp_data[1814] = 32'h522f2ab7;
temp_data[1815] = 32'h5237a9b5;
temp_data[1816] = 32'h52412168;
temp_data[1817] = 32'h524ba85d;
temp_data[1818] = 32'h525757ef;
temp_data[1819] = 32'h52644ca9;
temp_data[1820] = 32'h5272a687;
temp_data[1821] = 32'h52828955;
temp_data[1822] = 32'h52941d04;
temp_data[1823] = 32'h52a78e19;
temp_data[1824] = 32'h52bd0e2c;
temp_data[1825] = 32'h52d4d456;
temp_data[1826] = 32'h52ef1dd6;
temp_data[1827] = 32'h530c2e99;
temp_data[1828] = 32'h532c51f0;
temp_data[1829] = 32'h534fdb55;
temp_data[1830] = 32'h53772728;
temp_data[1831] = 32'h53a29baa;
temp_data[1832] = 32'h53d2a9e7;
temp_data[1833] = 32'h5407cf25;
temp_data[1834] = 32'h543e022a;
temp_data[1835] = 32'h546ef28c;
temp_data[1836] = 32'h549b202e;
temp_data[1837] = 32'h54c2fe5d;
temp_data[1838] = 32'h54e6f556;
temp_data[1839] = 32'h55076349;
temp_data[1840] = 32'h55249d49;
temp_data[1841] = 32'h553ef00b;
temp_data[1842] = 32'h5556a0c3;
temp_data[1843] = 32'h556bedc4;
temp_data[1844] = 32'h557f0f1f;
temp_data[1845] = 32'h55903733;
temp_data[1846] = 32'h559f9336;
temp_data[1847] = 32'h55ad4bad;
temp_data[1848] = 32'h55b984d3;
temp_data[1849] = 32'h55c45eee;
temp_data[1850] = 32'h55cdf6c7;
temp_data[1851] = 32'h55d665dc;
temp_data[1852] = 32'h55ddc2b1;
temp_data[1853] = 32'h55e4210c;
temp_data[1854] = 32'h55e99229;
temp_data[1855] = 32'h55ee24fb;
temp_data[1856] = 32'h55f1e636;
temp_data[1857] = 32'h55f4e09c;
temp_data[1858] = 32'h55f71cef;
temp_data[1859] = 32'h55f8a234;
temp_data[1860] = 32'h55f9759f;
temp_data[1861] = 32'h55f99acc;
temp_data[1862] = 32'h55f913a1;
temp_data[1863] = 32'h55f7e076;
temp_data[1864] = 32'h55f5fff8;
temp_data[1865] = 32'h55f36f3b;
temp_data[1866] = 32'h55f029aa;
temp_data[1867] = 32'h55ec28fe;
temp_data[1868] = 32'h55e76523;
temp_data[1869] = 32'h55e1d435;
temp_data[1870] = 32'h55db6a44;
temp_data[1871] = 32'h55d41954;
temp_data[1872] = 32'h55cbd12d;
temp_data[1873] = 32'h55c27f13;
temp_data[1874] = 32'h55b80dbf;
temp_data[1875] = 32'h55ac6502;
temp_data[1876] = 32'h559f698c;
temp_data[1877] = 32'h5590fca8;
temp_data[1878] = 32'h5580fbe3;
temp_data[1879] = 32'h556f40ab;
temp_data[1880] = 32'h555b9fe8;
temp_data[1881] = 32'h5545e996;
temp_data[1882] = 32'h552de83a;
temp_data[1883] = 32'h55136052;
temp_data[1884] = 32'h54f60fd0;
temp_data[1885] = 32'h54d5ad5c;
temp_data[1886] = 32'h54b1e7a3;
temp_data[1887] = 32'h548a6484;
temp_data[1888] = 32'h545ec040;
temp_data[1889] = 32'h542e8c69;
temp_data[1890] = 32'h53f94edb;
temp_data[1891] = 32'h53be800a;
temp_data[1892] = 32'h53870ae1;
temp_data[1893] = 32'h5354c250;
temp_data[1894] = 32'h532726e5;
temp_data[1895] = 32'h52fdc569;
temp_data[1896] = 32'h52d83598;
temp_data[1897] = 32'h52b6192f;
temp_data[1898] = 32'h52971ae7;
temp_data[1899] = 32'h527aedaf;
temp_data[1900] = 32'h52614be0;
temp_data[1901] = 32'h5249f690;
temp_data[1902] = 32'h5234b4fe;
temp_data[1903] = 32'h522153da;
temp_data[1904] = 32'h520fa4ec;
temp_data[1905] = 32'h51ff7e6f;
temp_data[1906] = 32'h51f0babf;
temp_data[1907] = 32'h51e337ef;
temp_data[1908] = 32'h51d6d75a;
temp_data[1909] = 32'h51cb7d6b;
temp_data[1910] = 32'h51c11141;
temp_data[1911] = 32'h51b77c63;
temp_data[1912] = 32'h51aeaa97;
temp_data[1913] = 32'h51a689a0;
temp_data[1914] = 32'h519f090b;
temp_data[1915] = 32'h519819fc;
temp_data[1916] = 32'h5191af0c;
temp_data[1917] = 32'h518bbc2c;
temp_data[1918] = 32'h5186366d;
temp_data[1919] = 32'h518113f9;
temp_data[1920] = 32'h517c4bec;
temp_data[1921] = 32'h5177d639;
temp_data[1922] = 32'h5173ab9f;
temp_data[1923] = 32'h516fc58b;
temp_data[1924] = 32'h516c1e11;
temp_data[1925] = 32'h5168afd1;
temp_data[1926] = 32'h516575ea;
temp_data[1927] = 32'h51626bfd;
temp_data[1928] = 32'h515f8e00;
temp_data[1929] = 32'h515cd862;
temp_data[1930] = 32'h515a47d0;
temp_data[1931] = 32'h5157d955;
temp_data[1932] = 32'h51558a3b;
temp_data[1933] = 32'h5153580c;
temp_data[1934] = 32'h5151408e;
temp_data[1935] = 32'h514f41b7;
temp_data[1936] = 32'h514d59b0;
temp_data[1937] = 32'h514b86c6;
temp_data[1938] = 32'h5149c76d;
temp_data[1939] = 32'h51481a3f;
temp_data[1940] = 32'h51467df6;
temp_data[1941] = 32'h5144f163;
temp_data[1942] = 32'h51437371;
temp_data[1943] = 32'h5142032e;
temp_data[1944] = 32'h51409fa5;
temp_data[1945] = 32'h513f480a;
temp_data[1946] = 32'h513dfb9c;
temp_data[1947] = 32'h513cb9a6;
temp_data[1948] = 32'h513b8184;
temp_data[1949] = 32'h513a529c;
temp_data[1950] = 32'h51392c62;
temp_data[1951] = 32'h51380e56;
temp_data[1952] = 32'h5136f7fd;
temp_data[1953] = 32'h5135e8ee;
temp_data[1954] = 32'h5134e0c1;
temp_data[1955] = 32'h5133df11;
temp_data[1956] = 32'h5132e38a;
temp_data[1957] = 32'h5131eddd;
temp_data[1958] = 32'h5130fdb5;
temp_data[1959] = 32'h513012cf;
temp_data[1960] = 32'h512f2ce9;
temp_data[1961] = 32'h512e4bc2;
temp_data[1962] = 32'h512d6f22;
temp_data[1963] = 32'h512c96d1;
temp_data[1964] = 32'h512bc29c;
temp_data[1965] = 32'h512af24e;
temp_data[1966] = 32'h512a25c0;
temp_data[1967] = 32'h51295cc0;
temp_data[1968] = 32'h5128972d;
temp_data[1969] = 32'h5127d4dc;
temp_data[1970] = 32'h512715ad;
temp_data[1971] = 32'h51265979;
temp_data[1972] = 32'h5125a01f;
temp_data[1973] = 32'h5124e985;
temp_data[1974] = 32'h5124358b;
temp_data[1975] = 32'h51238416;
temp_data[1976] = 32'h5122d50f;
temp_data[1977] = 32'h51222852;
temp_data[1978] = 32'h51217dd4;
temp_data[1979] = 32'h5120d573;
temp_data[1980] = 32'h51202f1f;
temp_data[1981] = 32'h511f8ac6;
temp_data[1982] = 32'h511ee84b;
temp_data[1983] = 32'h511e47a1;
temp_data[1984] = 32'h511da8b9;
temp_data[1985] = 32'h511d0b78;
temp_data[1986] = 32'h511c6fd2;
temp_data[1987] = 32'h511bd5bb;
temp_data[1988] = 32'h511b3d1d;
temp_data[1989] = 32'h511aa5ec;
temp_data[1990] = 32'h511a1017;
temp_data[1991] = 32'h51197b96;
temp_data[1992] = 32'h5118e857;
temp_data[1993] = 32'h5118564b;
temp_data[1994] = 32'h5117c56d;
temp_data[1995] = 32'h511735b1;
temp_data[1996] = 32'h5116a705;
temp_data[1997] = 32'h51161965;
temp_data[1998] = 32'h51158cc5;
temp_data[1999] = 32'h51150119;
temp_data[2000] = 32'h5114765c;
temp_data[2001] = 32'h5113ec85;
temp_data[2002] = 32'h51136388;
temp_data[2003] = 32'h5112db62;
temp_data[2004] = 32'h5112540d;
temp_data[2005] = 32'h5111cd7d;
temp_data[2006] = 32'h511147b6;
temp_data[2007] = 32'h5110c2a9;
temp_data[2008] = 32'h51103e57;
temp_data[2009] = 32'h510fbabf;
temp_data[2010] = 32'h510f37da;
temp_data[2011] = 32'h510eb5a6;
temp_data[2012] = 32'h510e3426;
temp_data[2013] = 32'h510db357;
temp_data[2014] = 32'h510d3340;
temp_data[2015] = 32'h510cb3dd;
temp_data[2016] = 32'h510c3533;
temp_data[2017] = 32'h510bb74e;
temp_data[2018] = 32'h510b3a2a;
temp_data[2019] = 32'h510abddc;
temp_data[2020] = 32'h510a4268;
temp_data[2021] = 32'h5109c7da;
temp_data[2022] = 32'h51094e40;
temp_data[2023] = 32'h5108d5b7;
temp_data[2024] = 32'h51085e46;
temp_data[2025] = 32'h5107e80c;
temp_data[2026] = 32'h51077326;
temp_data[2027] = 32'h5106ffb5;
temp_data[2028] = 32'h51068dd2;
temp_data[2029] = 32'h51061db4;
temp_data[2030] = 32'h5105af7d;
temp_data[2031] = 32'h5105436c;
temp_data[2032] = 32'h5104d9b2;
temp_data[2033] = 32'h51047297;
temp_data[2034] = 32'h51040e63;
temp_data[2035] = 32'h5103ad6d;
temp_data[2036] = 32'h5103500d;
temp_data[2037] = 32'h5102f6ad;
temp_data[2038] = 32'h5102a1c2;
temp_data[2039] = 32'h510251ce;
temp_data[2040] = 32'h51020768;
temp_data[2041] = 32'h5101c32b;
temp_data[2042] = 32'h510185cf;
temp_data[2043] = 32'h5101501e;
temp_data[2044] = 32'h510122fb;
temp_data[2045] = 32'h5100ff65;
temp_data[2046] = 32'h5100e671;
temp_data[2047] = 32'h5100d955;
temp_data[2048] = 32'h50f7069e;
temp_data[2049] = 32'h50f712f1;
temp_data[2050] = 32'h50f72a5e;
temp_data[2051] = 32'h50f74bb6;
temp_data[2052] = 32'h50f775e2;
temp_data[2053] = 32'h50f7a7eb;
temp_data[2054] = 32'h50f7e0f4;
temp_data[2055] = 32'h50f8203a;
temp_data[2056] = 32'h50f86506;
temp_data[2057] = 32'h50f8aebc;
temp_data[2058] = 32'h50f8fcce;
temp_data[2059] = 32'h50f94eba;
temp_data[2060] = 32'h50f9a40e;
temp_data[2061] = 32'h50f9fc65;
temp_data[2062] = 32'h50fa5764;
temp_data[2063] = 32'h50fab4b7;
temp_data[2064] = 32'h50fb1416;
temp_data[2065] = 32'h50fb7543;
temp_data[2066] = 32'h50fbd7fe;
temp_data[2067] = 32'h50fc3c19;
temp_data[2068] = 32'h50fca166;
temp_data[2069] = 32'h50fd07b8;
temp_data[2070] = 32'h50fd6eeb;
temp_data[2071] = 32'h50fdd6e0;
temp_data[2072] = 32'h50fe3f7d;
temp_data[2073] = 32'h50fea8a8;
temp_data[2074] = 32'h50ff124d;
temp_data[2075] = 32'h50ff7c52;
temp_data[2076] = 32'h50ffe6ac;
temp_data[2077] = 32'h51005148;
temp_data[2078] = 32'h5100bc1f;
temp_data[2079] = 32'h51012720;
temp_data[2080] = 32'h51019243;
temp_data[2081] = 32'h5101fd82;
temp_data[2082] = 32'h510268d7;
temp_data[2083] = 32'h5102d43d;
temp_data[2084] = 32'h51033fab;
temp_data[2085] = 32'h5103ab22;
temp_data[2086] = 32'h51041698;
temp_data[2087] = 32'h51048213;
temp_data[2088] = 32'h5104ed8d;
temp_data[2089] = 32'h51055908;
temp_data[2090] = 32'h5105c482;
temp_data[2091] = 32'h51062ff9;
temp_data[2092] = 32'h51069b74;
temp_data[2093] = 32'h510706ea;
temp_data[2094] = 32'h51077269;
temp_data[2095] = 32'h5107dde8;
temp_data[2096] = 32'h5108496f;
temp_data[2097] = 32'h5108b4fa;
temp_data[2098] = 32'h51092092;
temp_data[2099] = 32'h51098c37;
temp_data[2100] = 32'h5109f7ec;
temp_data[2101] = 32'h510a63b7;
temp_data[2102] = 32'h510acf96;
temp_data[2103] = 32'h510b3b8a;
temp_data[2104] = 32'h510ba7a0;
temp_data[2105] = 32'h510c13d3;
temp_data[2106] = 32'h510c802c;
temp_data[2107] = 32'h510cecab;
temp_data[2108] = 32'h510d5958;
temp_data[2109] = 32'h510dc632;
temp_data[2110] = 32'h510e3340;
temp_data[2111] = 32'h510ea084;
temp_data[2112] = 32'h510f0e06;
temp_data[2113] = 32'h510f7bc4;
temp_data[2114] = 32'h510fe9c9;
temp_data[2115] = 32'h51105819;
temp_data[2116] = 32'h5110c6b5;
temp_data[2117] = 32'h511135a0;
temp_data[2118] = 32'h5111a4e3;
temp_data[2119] = 32'h5112147f;
temp_data[2120] = 32'h5112847f;
temp_data[2121] = 32'h5112f4e0;
temp_data[2122] = 32'h511365ae;
temp_data[2123] = 32'h5113d6e9;
temp_data[2124] = 32'h51144899;
temp_data[2125] = 32'h5114bac3;
temp_data[2126] = 32'h51152d6b;
temp_data[2127] = 32'h5115a099;
temp_data[2128] = 32'h51161451;
temp_data[2129] = 32'h51168898;
temp_data[2130] = 32'h5116fd72;
temp_data[2131] = 32'h511772eb;
temp_data[2132] = 32'h5117e908;
temp_data[2133] = 32'h51185fc8;
temp_data[2134] = 32'h5118d73d;
temp_data[2135] = 32'h51194f61;
temp_data[2136] = 32'h5119c847;
temp_data[2137] = 32'h511a41f2;
temp_data[2138] = 32'h511abc62;
temp_data[2139] = 32'h511b37a8;
temp_data[2140] = 32'h511bb3cc;
temp_data[2141] = 32'h511c30cf;
temp_data[2142] = 32'h511caebc;
temp_data[2143] = 32'h511d2d9d;
temp_data[2144] = 32'h511dad7d;
temp_data[2145] = 32'h511e2e62;
temp_data[2146] = 32'h511eb057;
temp_data[2147] = 32'h511f336a;
temp_data[2148] = 32'h511fb79e;
temp_data[2149] = 32'h51203cff;
temp_data[2150] = 32'h5120c3a0;
temp_data[2151] = 32'h51214b84;
temp_data[2152] = 32'h5121d4bf;
temp_data[2153] = 32'h51225f5b;
temp_data[2154] = 32'h5122eb64;
temp_data[2155] = 32'h512378ea;
temp_data[2156] = 32'h512407fb;
temp_data[2157] = 32'h512498ab;
temp_data[2158] = 32'h51252b06;
temp_data[2159] = 32'h5125bf1f;
temp_data[2160] = 32'h51265508;
temp_data[2161] = 32'h5126ecd5;
temp_data[2162] = 32'h51278694;
temp_data[2163] = 32'h51282264;
temp_data[2164] = 32'h5128c055;
temp_data[2165] = 32'h51296080;
temp_data[2166] = 32'h512a02fb;
temp_data[2167] = 32'h512aa7e3;
temp_data[2168] = 32'h512b4f4c;
temp_data[2169] = 32'h512bf959;
temp_data[2170] = 32'h512ca622;
temp_data[2171] = 32'h512d55c5;
temp_data[2172] = 32'h512e0863;
temp_data[2173] = 32'h512ebe16;
temp_data[2174] = 32'h512f7708;
temp_data[2175] = 32'h51303351;
temp_data[2176] = 32'h5130f317;
temp_data[2177] = 32'h5131b680;
temp_data[2178] = 32'h51327daa;
temp_data[2179] = 32'h513348b6;
temp_data[2180] = 32'h513417ce;
temp_data[2181] = 32'h5134eb10;
temp_data[2182] = 32'h5135c298;
temp_data[2183] = 32'h51369e8c;
temp_data[2184] = 32'h51377f02;
temp_data[2185] = 32'h51386417;
temp_data[2186] = 32'h51394ddb;
temp_data[2187] = 32'h513a3c60;
temp_data[2188] = 32'h513b2fad;
temp_data[2189] = 32'h513c27c4;
temp_data[2190] = 32'h513d249e;
temp_data[2191] = 32'h513e2629;
temp_data[2192] = 32'h513f2c45;
temp_data[2193] = 32'h514036c6;
temp_data[2194] = 32'h51414574;
temp_data[2195] = 32'h51425800;
temp_data[2196] = 32'h51436e11;
temp_data[2197] = 32'h51448733;
temp_data[2198] = 32'h5145a2e0;
temp_data[2199] = 32'h5146c083;
temp_data[2200] = 32'h5147df6a;
temp_data[2201] = 32'h5148fed2;
temp_data[2202] = 32'h514a1deb;
temp_data[2203] = 32'h514b3bc5;
temp_data[2204] = 32'h514c576d;
temp_data[2205] = 32'h514d717a;
temp_data[2206] = 32'h514e8f58;
temp_data[2207] = 32'h514fb00c;
temp_data[2208] = 32'h5150d2a2;
temp_data[2209] = 32'h5151f640;
temp_data[2210] = 32'h51531a1e;
temp_data[2211] = 32'h51543d86;
temp_data[2212] = 32'h51555fdd;
temp_data[2213] = 32'h5156809d;
temp_data[2214] = 32'h51579f51;
temp_data[2215] = 32'h5158bba1;
temp_data[2216] = 32'h5159d545;
temp_data[2217] = 32'h515aec0b;
temp_data[2218] = 32'h515bffce;
temp_data[2219] = 32'h515d1084;
temp_data[2220] = 32'h515e1e26;
temp_data[2221] = 32'h515f28c3;
temp_data[2222] = 32'h5160307b;
temp_data[2223] = 32'h5161356e;
temp_data[2224] = 32'h516237ca;
temp_data[2225] = 32'h516337ce;
temp_data[2226] = 32'h516435b9;
temp_data[2227] = 32'h516531db;
temp_data[2228] = 32'h51662c84;
temp_data[2229] = 32'h5167260f;
temp_data[2230] = 32'h51681ee2;
temp_data[2231] = 32'h5169176a;
temp_data[2232] = 32'h516a1017;
temp_data[2233] = 32'h516b0963;
temp_data[2234] = 32'h516c03da;
temp_data[2235] = 32'h516d0004;
temp_data[2236] = 32'h516dfe82;
temp_data[2237] = 32'h516efff3;
temp_data[2238] = 32'h5170050c;
temp_data[2239] = 32'h51710e91;
temp_data[2240] = 32'h51721d54;
temp_data[2241] = 32'h51733233;
temp_data[2242] = 32'h51744e27;
temp_data[2243] = 32'h51757243;
temp_data[2244] = 32'h51769fa9;
temp_data[2245] = 32'h5177d799;
temp_data[2246] = 32'h51791b7a;
temp_data[2247] = 32'h517a6cce;
temp_data[2248] = 32'h517bcd3e;
temp_data[2249] = 32'h517d3e9f;
temp_data[2250] = 32'h517ec2fc;
temp_data[2251] = 32'h51805c8e;
temp_data[2252] = 32'h51820dcc;
temp_data[2253] = 32'h5183d96a;
temp_data[2254] = 32'h5185c276;
temp_data[2255] = 32'h5187cc42;
temp_data[2256] = 32'h5189fa7f;
temp_data[2257] = 32'h518c5144;
temp_data[2258] = 32'h518ed51b;
temp_data[2259] = 32'h51918b0d;
temp_data[2260] = 32'h519478ab;
temp_data[2261] = 32'h5197a427;
temp_data[2262] = 32'h519b1455;
temp_data[2263] = 32'h519ed0d9;
temp_data[2264] = 32'h51a2e219;
temp_data[2265] = 32'h51a7516e;
temp_data[2266] = 32'h51ac292c;
temp_data[2267] = 32'h51b174d1;
temp_data[2268] = 32'h51b74107;
temp_data[2269] = 32'h51bd9bdc;
temp_data[2270] = 32'h51c494d9;
temp_data[2271] = 32'h51cc3d29;
temp_data[2272] = 32'h51d4a7c6;
temp_data[2273] = 32'h51dde99f;
temp_data[2274] = 32'h51e819db;
temp_data[2275] = 32'h51f35215;
temp_data[2276] = 32'h51fdd790;
temp_data[2277] = 32'h52074ef9;
temp_data[2278] = 32'h520fcfff;
temp_data[2279] = 32'h52176fb5;
temp_data[2280] = 32'h521e40ea;
temp_data[2281] = 32'h52245443;
temp_data[2282] = 32'h5229b86f;
temp_data[2283] = 32'h522e7a42;
temp_data[2284] = 32'h5232a4d7;
temp_data[2285] = 32'h523641af;
temp_data[2286] = 32'h523958c9;
temp_data[2287] = 32'h523bf0b3;
temp_data[2288] = 32'h523e0ea2;
temp_data[2289] = 32'h523fb670;
temp_data[2290] = 32'h5240eabc;
temp_data[2291] = 32'h5241aceb;
temp_data[2292] = 32'h5241fd2a;
temp_data[2293] = 32'h5241da66;
temp_data[2294] = 32'h52414268;
temp_data[2295] = 32'h524031a9;
temp_data[2296] = 32'h523ea372;
temp_data[2297] = 32'h523c91b0;
temp_data[2298] = 32'h5239f4fd;
temp_data[2299] = 32'h5236c482;
temp_data[2300] = 32'h5232f5e8;
temp_data[2301] = 32'h522e7d31;
temp_data[2302] = 32'h52294cad;
temp_data[2303] = 32'h522354ca;
temp_data[2304] = 32'h521c83d8;
temp_data[2305] = 32'h52169b89;
temp_data[2306] = 32'h52118a4c;
temp_data[2307] = 32'h520d40b8;
temp_data[2308] = 32'h5209b16c;
temp_data[2309] = 32'h5206d0cc;
temp_data[2310] = 32'h52049503;
temp_data[2311] = 32'h5202f5d3;
temp_data[2312] = 32'h5201ec89;
temp_data[2313] = 32'h520173f3;
temp_data[2314] = 32'h52018848;
temp_data[2315] = 32'h5202272d;
temp_data[2316] = 32'h52034fa5;
temp_data[2317] = 32'h5205020c;
temp_data[2318] = 32'h52074035;
temp_data[2319] = 32'h520a0d4e;
temp_data[2320] = 32'h520d6e01;
temp_data[2321] = 32'h52116877;
temp_data[2322] = 32'h52160475;
temp_data[2323] = 32'h521b4b62;
temp_data[2324] = 32'h5221487c;
temp_data[2325] = 32'h522808dd;
temp_data[2326] = 32'h522f9bb2;
temp_data[2327] = 32'h5238125e;
temp_data[2328] = 32'h524180b2;
temp_data[2329] = 32'h524bfd1a;
temp_data[2330] = 32'h5257a0f1;
temp_data[2331] = 32'h526488a4;
temp_data[2332] = 32'h5272d428;
temp_data[2333] = 32'h5282a733;
temp_data[2334] = 32'h529429ae;
temp_data[2335] = 32'h52a7881a;
temp_data[2336] = 32'h52bcf402;
temp_data[2337] = 32'h52d4a490;
temp_data[2338] = 32'h52eed6fe;
temp_data[2339] = 32'h530bcf57;
temp_data[2340] = 32'h532bd902;
temp_data[2341] = 32'h534f4795;
temp_data[2342] = 32'h537677a3;
temp_data[2343] = 32'h53a1cf9a;
temp_data[2344] = 32'h53d1c0c2;
temp_data[2345] = 32'h5406c897;
temp_data[2346] = 32'h543cde22;
temp_data[2347] = 32'h546db142;
temp_data[2348] = 32'h5499c20d;
temp_data[2349] = 32'h54c1840e;
temp_data[2350] = 32'h54e55fb3;
temp_data[2351] = 32'h5505b35b;
temp_data[2352] = 32'h5522d439;
temp_data[2353] = 32'h553d0f1f;
temp_data[2354] = 32'h5554a958;
temp_data[2355] = 32'h5569e13f;
temp_data[2356] = 32'h557ceeee;
temp_data[2357] = 32'h558e04bc;
temp_data[2358] = 32'h559d4fdf;
temp_data[2359] = 32'h55aaf8d3;
temp_data[2360] = 32'h55b723bc;
temp_data[2361] = 32'h55c1f0e1;
temp_data[2362] = 32'h55cb7cf2;
temp_data[2363] = 32'h55d3e15d;
temp_data[2364] = 32'h55db3498;
temp_data[2365] = 32'h55e18a55;
temp_data[2366] = 32'h55e6f3cb;
temp_data[2367] = 32'h55eb7fd8;
temp_data[2368] = 32'h55ef3b2a;
temp_data[2369] = 32'h55f2306a;
temp_data[2370] = 32'h55f4685e;
temp_data[2371] = 32'h55f5e9fb;
temp_data[2372] = 32'h55f6ba77;
temp_data[2373] = 32'h55f6dd61;
temp_data[2374] = 32'h55f654a0;
temp_data[2375] = 32'h55f52086;
temp_data[2376] = 32'h55f33fc8;
temp_data[2377] = 32'h55f0af75;
temp_data[2378] = 32'h55ed6b05;
temp_data[2379] = 32'h55e96c2b;
temp_data[2380] = 32'h55e4aae7;
temp_data[2381] = 32'h55df1d50;
temp_data[2382] = 32'h55d8b78d;
temp_data[2383] = 32'h55d16ba5;
temp_data[2384] = 32'h55c9296f;
temp_data[2385] = 32'h55bfde44;
temp_data[2386] = 32'h55b574eb;
temp_data[2387] = 32'h55a9d539;
temp_data[2388] = 32'h559ce400;
temp_data[2389] = 32'h558e828c;
temp_data[2390] = 32'h557e8e7e;
temp_data[2391] = 32'h556ce150;
temp_data[2392] = 32'h55594ff4;
temp_data[2393] = 32'h5543aa6d;
temp_data[2394] = 32'h552bbb3d;
temp_data[2395] = 32'h551146e5;
temp_data[2396] = 32'h54f40b46;
temp_data[2397] = 32'h54d3bef5;
temp_data[2398] = 32'h54b01080;
temp_data[2399] = 32'h5488a5a9;
temp_data[2400] = 32'h545d1a82;
temp_data[2401] = 32'h542d006d;
temp_data[2402] = 32'h53f7dd09;
temp_data[2403] = 32'h53bd2895;
temp_data[2404] = 32'h5385cdb8;
temp_data[2405] = 32'h53539f27;
temp_data[2406] = 32'h53261d36;
temp_data[2407] = 32'h52fcd478;
temp_data[2408] = 32'h52d75c81;
temp_data[2409] = 32'h52b556e2;
temp_data[2410] = 32'h52966e37;
temp_data[2411] = 32'h527a5554;
temp_data[2412] = 32'h5260c68f;
temp_data[2413] = 32'h524982f5;
temp_data[2414] = 32'h523451bd;
temp_data[2415] = 32'h5220ffa8;
temp_data[2416] = 32'h520f5e7d;
temp_data[2417] = 32'h51ff4489;
temp_data[2418] = 32'h51f08c3b;
temp_data[2419] = 32'h51e313b2;
temp_data[2420] = 32'h51d6bc62;
temp_data[2421] = 32'h51cb6abe;
temp_data[2422] = 32'h51c105ff;
temp_data[2423] = 32'h51b777c0;
temp_data[2424] = 32'h51aeabd6;
temp_data[2425] = 32'h51a69015;
temp_data[2426] = 32'h519f1416;
temp_data[2427] = 32'h51982913;
temp_data[2428] = 32'h5191c1b1;
temp_data[2429] = 32'h518bd1e5;
temp_data[2430] = 32'h51864edb;
temp_data[2431] = 32'h51812eba;
temp_data[2432] = 32'h517c68ad;
temp_data[2433] = 32'h5177f4b2;
temp_data[2434] = 32'h5173cb8e;
temp_data[2435] = 32'h516fe6b8;
temp_data[2436] = 32'h516c4042;
temp_data[2437] = 32'h5168d2d8;
temp_data[2438] = 32'h516599a2;
temp_data[2439] = 32'h5162903a;
temp_data[2440] = 32'h515fb2ab;
temp_data[2441] = 32'h515cfd54;
temp_data[2442] = 32'h515a6cf4;
temp_data[2443] = 32'h5157fe97;
temp_data[2444] = 32'h5155af86;
temp_data[2445] = 32'h51537d4e;
temp_data[2446] = 32'h515165b6;
temp_data[2447] = 32'h514f66ba;
temp_data[2448] = 32'h514d7e80;
temp_data[2449] = 32'h514bab54;
temp_data[2450] = 32'h5149ebb7;
temp_data[2451] = 32'h51483e3e;
temp_data[2452] = 32'h5146a19d;
temp_data[2453] = 32'h514514b1;
temp_data[2454] = 32'h51439664;
temp_data[2455] = 32'h514225b7;
temp_data[2456] = 32'h5140c1c6;
temp_data[2457] = 32'h513f69c2;
temp_data[2458] = 32'h513e1ce7;
temp_data[2459] = 32'h513cda7f;
temp_data[2460] = 32'h513ba1ec;
temp_data[2461] = 32'h513a728f;
temp_data[2462] = 32'h51394be0;
temp_data[2463] = 32'h51382d5e;
temp_data[2464] = 32'h51371694;
temp_data[2465] = 32'h5136070c;
temp_data[2466] = 32'h5134fe65;
temp_data[2467] = 32'h5133fc44;
temp_data[2468] = 32'h51330047;
temp_data[2469] = 32'h51320a20;
temp_data[2470] = 32'h51311983;
temp_data[2471] = 32'h51302e27;
temp_data[2472] = 32'h512f47cb;
temp_data[2473] = 32'h512e6630;
temp_data[2474] = 32'h512d891a;
temp_data[2475] = 32'h512cb053;
temp_data[2476] = 32'h512bdba9;
temp_data[2477] = 32'h512b0ae9;
temp_data[2478] = 32'h512a3dea;
temp_data[2479] = 32'h51297479;
temp_data[2480] = 32'h5128ae75;
temp_data[2481] = 32'h5127ebb7;
temp_data[2482] = 32'h51272c17;
temp_data[2483] = 32'h51266f72;
temp_data[2484] = 32'h5125b5af;
temp_data[2485] = 32'h5124fea8;
temp_data[2486] = 32'h51244a41;
temp_data[2487] = 32'h51239863;
temp_data[2488] = 32'h5122e8ee;
temp_data[2489] = 32'h51223bc9;
temp_data[2490] = 32'h512190de;
temp_data[2491] = 32'h5120e819;
temp_data[2492] = 32'h5120415f;
temp_data[2493] = 32'h511f9c9d;
temp_data[2494] = 32'h511ef9be;
temp_data[2495] = 32'h511e58b0;
temp_data[2496] = 32'h511db963;
temp_data[2497] = 32'h511d1bbd;
temp_data[2498] = 32'h511c7fb7;
temp_data[2499] = 32'h511be53b;
temp_data[2500] = 32'h511b4c3c;
temp_data[2501] = 32'h511ab4ab;
temp_data[2502] = 32'h511a1e75;
temp_data[2503] = 32'h51198994;
temp_data[2504] = 32'h5118f5f5;
temp_data[2505] = 32'h51186391;
temp_data[2506] = 32'h5117d252;
temp_data[2507] = 32'h51174239;
temp_data[2508] = 32'h5116b331;
temp_data[2509] = 32'h51162535;
temp_data[2510] = 32'h51159839;
temp_data[2511] = 32'h51150c35;
temp_data[2512] = 32'h5114811f;
temp_data[2513] = 32'h5113f6ec;
temp_data[2514] = 32'h51136d98;
temp_data[2515] = 32'h5112e519;
temp_data[2516] = 32'h51125d6c;
temp_data[2517] = 32'h5111d688;
temp_data[2518] = 32'h5111506a;
temp_data[2519] = 32'h5110cb08;
temp_data[2520] = 32'h5110465f;
temp_data[2521] = 32'h510fc272;
temp_data[2522] = 32'h510f3f3a;
temp_data[2523] = 32'h510ebcb2;
temp_data[2524] = 32'h510e3ae2;
temp_data[2525] = 32'h510db9bf;
temp_data[2526] = 32'h510d3954;
temp_data[2527] = 32'h510cb9a1;
temp_data[2528] = 32'h510c3aac;
temp_data[2529] = 32'h510bbc73;
temp_data[2530] = 32'h510b3f03;
temp_data[2531] = 32'h510ac265;
temp_data[2532] = 32'h510a46a2;
temp_data[2533] = 32'h5109cbc9;
temp_data[2534] = 32'h510951e7;
temp_data[2535] = 32'h5108d90e;
temp_data[2536] = 32'h51086156;
temp_data[2537] = 32'h5107ead5;
temp_data[2538] = 32'h510775a7;
temp_data[2539] = 32'h510701eb;
temp_data[2540] = 32'h51068fc9;
temp_data[2541] = 32'h51061f64;
temp_data[2542] = 32'h5105b0ee;
temp_data[2543] = 32'h5105449a;
temp_data[2544] = 32'h5104daa1;
temp_data[2545] = 32'h51047347;
temp_data[2546] = 32'h51040edc;
temp_data[2547] = 32'h5103adac;
temp_data[2548] = 32'h51035012;
temp_data[2549] = 32'h5102f67f;
temp_data[2550] = 32'h5102a162;
temp_data[2551] = 32'h51025144;
temp_data[2552] = 32'h510206af;
temp_data[2553] = 32'h5101c24c;
temp_data[2554] = 32'h510184cf;
temp_data[2555] = 32'h51014f01;
temp_data[2556] = 32'h510121c4;
temp_data[2557] = 32'h5100fe1e;
temp_data[2558] = 32'h5100e51d;
temp_data[2559] = 32'h5100d7fe;
temp_data[2560] = 32'h50f6fda0;
temp_data[2561] = 32'h50f709f6;
temp_data[2562] = 32'h50f7216c;
temp_data[2563] = 32'h50f742d5;
temp_data[2564] = 32'h50f76d11;
temp_data[2565] = 32'h50f79f38;
temp_data[2566] = 32'h50f7d862;
temp_data[2567] = 32'h50f817c6;
temp_data[2568] = 32'h50f85cbc;
temp_data[2569] = 32'h50f8a69c;
temp_data[2570] = 32'h50f8f4dc;
temp_data[2571] = 32'h50f946fa;
temp_data[2572] = 32'h50f99c84;
temp_data[2573] = 32'h50f9f512;
temp_data[2574] = 32'h50fa504c;
temp_data[2575] = 32'h50faadda;
temp_data[2576] = 32'h50fb0d78;
temp_data[2577] = 32'h50fb6ee3;
temp_data[2578] = 32'h50fbd1e1;
temp_data[2579] = 32'h50fc363f;
temp_data[2580] = 32'h50fc9bd0;
temp_data[2581] = 32'h50fd0269;
temp_data[2582] = 32'h50fd69e4;
temp_data[2583] = 32'h50fdd224;
temp_data[2584] = 32'h50fe3b08;
temp_data[2585] = 32'h50fea47f;
temp_data[2586] = 32'h50ff0e6b;
temp_data[2587] = 32'h50ff78c0;
temp_data[2588] = 32'h50ffe365;
temp_data[2589] = 32'h51004e51;
temp_data[2590] = 32'h5100b973;
temp_data[2591] = 32'h510124c4;
temp_data[2592] = 32'h5101903a;
temp_data[2593] = 32'h5101fbca;
temp_data[2594] = 32'h51026773;
temp_data[2595] = 32'h5102d328;
temp_data[2596] = 32'h51033ee6;
temp_data[2597] = 32'h5103aab0;
temp_data[2598] = 32'h5104167b;
temp_data[2599] = 32'h51048249;
temp_data[2600] = 32'h5104ee18;
temp_data[2601] = 32'h510559e6;
temp_data[2602] = 32'h5105c5b5;
temp_data[2603] = 32'h51063183;
temp_data[2604] = 32'h51069d52;
temp_data[2605] = 32'h51070920;
temp_data[2606] = 32'h510774f3;
temp_data[2607] = 32'h5107e0ca;
temp_data[2608] = 32'h51084ca9;
temp_data[2609] = 32'h5108b88d;
temp_data[2610] = 32'h5109247d;
temp_data[2611] = 32'h5109907e;
temp_data[2612] = 32'h5109fc8b;
temp_data[2613] = 32'h510a68ad;
temp_data[2614] = 32'h510ad4e5;
temp_data[2615] = 32'h510b4135;
temp_data[2616] = 32'h510bada7;
temp_data[2617] = 32'h510c1a37;
temp_data[2618] = 32'h510c86e8;
temp_data[2619] = 32'h510cf3c7;
temp_data[2620] = 32'h510d60cc;
temp_data[2621] = 32'h510dce03;
temp_data[2622] = 32'h510e3b71;
temp_data[2623] = 32'h510ea915;
temp_data[2624] = 32'h510f16f4;
temp_data[2625] = 32'h510f8512;
temp_data[2626] = 32'h510ff377;
temp_data[2627] = 32'h51106224;
temp_data[2628] = 32'h5110d120;
temp_data[2629] = 32'h51114070;
temp_data[2630] = 32'h5111b014;
temp_data[2631] = 32'h51122014;
temp_data[2632] = 32'h51129075;
temp_data[2633] = 32'h5113013f;
temp_data[2634] = 32'h51137271;
temp_data[2635] = 32'h5113e411;
temp_data[2636] = 32'h5114562a;
temp_data[2637] = 32'h5114c8b8;
temp_data[2638] = 32'h51153bc9;
temp_data[2639] = 32'h5115af60;
temp_data[2640] = 32'h51162381;
temp_data[2641] = 32'h51169831;
temp_data[2642] = 32'h51170d78;
temp_data[2643] = 32'h5117835e;
temp_data[2644] = 32'h5117f9e8;
temp_data[2645] = 32'h51187119;
temp_data[2646] = 32'h5118e8fb;
temp_data[2647] = 32'h51196191;
temp_data[2648] = 32'h5119dae8;
temp_data[2649] = 32'h511a5504;
temp_data[2650] = 32'h511acfee;
temp_data[2651] = 32'h511b4ba9;
temp_data[2652] = 32'h511bc843;
temp_data[2653] = 32'h511c45bf;
temp_data[2654] = 32'h511cc426;
temp_data[2655] = 32'h511d4389;
temp_data[2656] = 32'h511dc3e3;
temp_data[2657] = 32'h511e454a;
temp_data[2658] = 32'h511ec7c1;
temp_data[2659] = 32'h511f4b55;
temp_data[2660] = 32'h511fd014;
temp_data[2661] = 32'h51205600;
temp_data[2662] = 32'h5120dd2b;
temp_data[2663] = 32'h512165a1;
temp_data[2664] = 32'h5121ef6b;
temp_data[2665] = 32'h51227a9e;
temp_data[2666] = 32'h5123073e;
temp_data[2667] = 32'h51239564;
temp_data[2668] = 32'h51242518;
temp_data[2669] = 32'h5124b66b;
temp_data[2670] = 32'h5125496f;
temp_data[2671] = 32'h5125de37;
temp_data[2672] = 32'h512674d6;
temp_data[2673] = 32'h51270d5f;
temp_data[2674] = 32'h5127a7e3;
temp_data[2675] = 32'h5128447c;
temp_data[2676] = 32'h5128e33f;
temp_data[2677] = 32'h51298445;
temp_data[2678] = 32'h512a27a6;
temp_data[2679] = 32'h512acd7d;
temp_data[2680] = 32'h512b75e2;
temp_data[2681] = 32'h512c20f7;
temp_data[2682] = 32'h512cced9;
temp_data[2683] = 32'h512d7fa2;
temp_data[2684] = 32'h512e3376;
temp_data[2685] = 32'h512eea79;
temp_data[2686] = 32'h512fa4ca;
temp_data[2687] = 32'h5130628d;
temp_data[2688] = 32'h513123e6;
temp_data[2689] = 32'h5131e8ff;
temp_data[2690] = 32'h5132b1fb;
temp_data[2691] = 32'h51337efe;
temp_data[2692] = 32'h5134502f;
temp_data[2693] = 32'h513525b3;
temp_data[2694] = 32'h5135ffb5;
temp_data[2695] = 32'h5136de51;
temp_data[2696] = 32'h5137c1a9;
temp_data[2697] = 32'h5138a9da;
temp_data[2698] = 32'h51399703;
temp_data[2699] = 32'h513a8937;
temp_data[2700] = 32'h513b8080;
temp_data[2701] = 32'h513c7cee;
temp_data[2702] = 32'h513d7e74;
temp_data[2703] = 32'h513e850e;
temp_data[2704] = 32'h513f909f;
temp_data[2705] = 32'h5140a101;
temp_data[2706] = 32'h5141b5fa;
temp_data[2707] = 32'h5142cf46;
temp_data[2708] = 32'h5143ec85;
temp_data[2709] = 32'h51450d45;
temp_data[2710] = 32'h514630fd;
temp_data[2711] = 32'h51475708;
temp_data[2712] = 32'h51487eb7;
temp_data[2713] = 32'h5149a72f;
temp_data[2714] = 32'h514acf96;
temp_data[2715] = 32'h514bf6ec;
temp_data[2716] = 32'h514d1c2e;
temp_data[2717] = 32'h514e3fd9;
temp_data[2718] = 32'h514f6745;
temp_data[2719] = 32'h51509160;
temp_data[2720] = 32'h5151bd2b;
temp_data[2721] = 32'h5152e9bc;
temp_data[2722] = 32'h51541633;
temp_data[2723] = 32'h515541d9;
temp_data[2724] = 32'h51566c05;
temp_data[2725] = 32'h51579429;
temp_data[2726] = 32'h5158b9d4;
temp_data[2727] = 32'h5159dca5;
temp_data[2728] = 32'h515afc59;
temp_data[2729] = 32'h515c18c2;
temp_data[2730] = 32'h515d31be;
temp_data[2731] = 32'h515e4741;
temp_data[2732] = 32'h515f5953;
temp_data[2733] = 32'h5160680a;
temp_data[2734] = 32'h5161737e;
temp_data[2735] = 32'h51627bdd;
temp_data[2736] = 32'h5163815a;
temp_data[2737] = 32'h5164843c;
temp_data[2738] = 32'h516584c7;
temp_data[2739] = 32'h5166834d;
temp_data[2740] = 32'h5167801f;
temp_data[2741] = 32'h51687ba6;
temp_data[2742] = 32'h51697647;
temp_data[2743] = 32'h516a7069;
temp_data[2744] = 32'h516b6a8c;
temp_data[2745] = 32'h516c652c;
temp_data[2746] = 32'h516d60cc;
temp_data[2747] = 32'h516e5e03;
temp_data[2748] = 32'h516f5d68;
temp_data[2749] = 32'h51705fa2;
temp_data[2750] = 32'h5171656b;
temp_data[2751] = 32'h51726f7a;
temp_data[2752] = 32'h51737eaa;
temp_data[2753] = 32'h517493de;
temp_data[2754] = 32'h5175b008;
temp_data[2755] = 32'h5176d435;
temp_data[2756] = 32'h5178018e;
temp_data[2757] = 32'h51793954;
temp_data[2758] = 32'h517a7ce5;
temp_data[2759] = 32'h517bcdc4;
temp_data[2760] = 32'h517d2d99;
temp_data[2761] = 32'h517e9e38;
temp_data[2762] = 32'h518021a3;
temp_data[2763] = 32'h5181ba13;
temp_data[2764] = 32'h518369fd;
temp_data[2765] = 32'h51853411;
temp_data[2766] = 32'h51871b58;
temp_data[2767] = 32'h5189231c;
temp_data[2768] = 32'h518b4f0e;
temp_data[2769] = 32'h518da340;
temp_data[2770] = 32'h51902435;
temp_data[2771] = 32'h5192d6ed;
temp_data[2772] = 32'h5195c0fd;
temp_data[2773] = 32'h5198e886;
temp_data[2774] = 32'h519c5469;
temp_data[2775] = 32'h51a00c31;
temp_data[2776] = 32'h51a41850;
temp_data[2777] = 32'h51a88217;
temp_data[2778] = 32'h51ad53e3;
temp_data[2779] = 32'h51b29928;
temp_data[2780] = 32'h51b85e9e;
temp_data[2781] = 32'h51beb257;
temp_data[2782] = 32'h51c5a3e8;
temp_data[2783] = 32'h51cd4480;
temp_data[2784] = 32'h51d5a733;
temp_data[2785] = 32'h51dee100;
temp_data[2786] = 32'h51e90920;
temp_data[2787] = 32'h51f43947;
temp_data[2788] = 32'h51feb6c8;
temp_data[2789] = 32'h5208266c;
temp_data[2790] = 32'h52109ff1;
temp_data[2791] = 32'h52183882;
temp_data[2792] = 32'h521f0300;
temp_data[2793] = 32'h5225101b;
temp_data[2794] = 32'h522a6e87;
temp_data[2795] = 32'h522f2b28;
temp_data[2796] = 32'h5233511a;
temp_data[2797] = 32'h5236e9e2;
temp_data[2798] = 32'h5239fd7e;
temp_data[2799] = 32'h523c9279;
temp_data[2800] = 32'h523eae00;
temp_data[2801] = 32'h524053f4;
temp_data[2802] = 32'h524186e8;
temp_data[2803] = 32'h52424834;
temp_data[2804] = 32'h52429803;
temp_data[2805] = 32'h5242753a;
temp_data[2806] = 32'h5241dd94;
temp_data[2807] = 32'h5240cd8e;
temp_data[2808] = 32'h523f4057;
temp_data[2809] = 32'h523d2fdc;
temp_data[2810] = 32'h523a94af;
temp_data[2811] = 32'h523765ed;
temp_data[2812] = 32'h52339935;
temp_data[2813] = 32'h522f2281;
temp_data[2814] = 32'h5229f417;
temp_data[2815] = 32'h5223fe58;
temp_data[2816] = 32'h521d2f8c;
temp_data[2817] = 32'h52174962;
temp_data[2818] = 32'h52123a36;
temp_data[2819] = 32'h520df29d;
temp_data[2820] = 32'h520a6523;
temp_data[2821] = 32'h52078627;
temp_data[2822] = 32'h52054bcb;
temp_data[2823] = 32'h5203adc1;
temp_data[2824] = 32'h5202a551;
temp_data[2825] = 32'h52022d3c;
temp_data[2826] = 32'h520241ab;
temp_data[2827] = 32'h5202e037;
temp_data[2828] = 32'h520407d5;
temp_data[2829] = 32'h5205b8dc;
temp_data[2830] = 32'h5207f50a;
temp_data[2831] = 32'h520abf7b;
temp_data[2832] = 32'h520e1cd2;
temp_data[2833] = 32'h5212131f;
temp_data[2834] = 32'h5216aa19;
temp_data[2835] = 32'h521beb18;
temp_data[2836] = 32'h5221e13b;
temp_data[2837] = 32'h52289991;
temp_data[2838] = 32'h5230232d;
temp_data[2839] = 32'h52388f60;
temp_data[2840] = 32'h5241f1d8;
temp_data[2841] = 32'h524c60fa;
temp_data[2842] = 32'h5257f5f5;
temp_data[2843] = 32'h5264cd31;
temp_data[2844] = 32'h52730681;
temp_data[2845] = 32'h5282c58f;
temp_data[2846] = 32'h5294322f;
temp_data[2847] = 32'h52a778dd;
temp_data[2848] = 32'h52bccb19;
temp_data[2849] = 32'h52d4600f;
temp_data[2850] = 32'h52ee750c;
temp_data[2851] = 32'h530b4e27;
temp_data[2852] = 32'h532b36eb;
temp_data[2853] = 32'h534e831f;
temp_data[2854] = 32'h53758f82;
temp_data[2855] = 32'h53a0c2ca;
temp_data[2856] = 32'h53d08e8a;
temp_data[2857] = 32'h5405708f;
temp_data[2858] = 32'h543b6035;
temp_data[2859] = 32'h546c0db2;
temp_data[2860] = 32'h5497f96e;
temp_data[2861] = 32'h54bf973e;
temp_data[2862] = 32'h54e34fdb;
temp_data[2863] = 32'h550381d4;
temp_data[2864] = 32'h55208290;
temp_data[2865] = 32'h553a9f06;
temp_data[2866] = 32'h55521c93;
temp_data[2867] = 32'h5567399f;
temp_data[2868] = 32'h557a2e49;
temp_data[2869] = 32'h558b2ced;
temp_data[2870] = 32'h559a62b2;
temp_data[2871] = 32'h55a7f7fd;
temp_data[2872] = 32'h55b410f1;
temp_data[2873] = 32'h55becdb8;
temp_data[2874] = 32'h55c84aed;
temp_data[2875] = 32'h55d0a1ec;
temp_data[2876] = 32'h55d7e914;
temp_data[2877] = 32'h55de3405;
temp_data[2878] = 32'h55e393e2;
temp_data[2879] = 32'h55e8176e;
temp_data[2880] = 32'h55ebcb4f;
temp_data[2881] = 32'h55eeba23;
temp_data[2882] = 32'h55f0eca2;
temp_data[2883] = 32'h55f269ad;
temp_data[2884] = 32'h55f3367e;
temp_data[2885] = 32'h55f35697;
temp_data[2886] = 32'h55f2cbde;
temp_data[2887] = 32'h55f196a2;
temp_data[2888] = 32'h55efb59a;
temp_data[2889] = 32'h55ed25d9;
temp_data[2890] = 32'h55e9e2d6;
temp_data[2891] = 32'h55e5e64f;
temp_data[2892] = 32'h55e1284e;
temp_data[2893] = 32'h55db9ef5;
temp_data[2894] = 32'h55d53e79;
temp_data[2895] = 32'h55cdf8f4;
temp_data[2896] = 32'h55c5be44;
temp_data[2897] = 32'h55bc7bdd;
temp_data[2898] = 32'h55b21c97;
temp_data[2899] = 32'h55a68861;
temp_data[2900] = 32'h5599a41a;
temp_data[2901] = 32'h558b512f;
temp_data[2902] = 32'h557b6d44;
temp_data[2903] = 32'h5569d1f2;
temp_data[2904] = 32'h55565437;
temp_data[2905] = 32'h5540c41a;
temp_data[2906] = 32'h5528ec25;
temp_data[2907] = 32'h550e90d1;
temp_data[2908] = 32'h54f16ff4;
temp_data[2909] = 32'h54d14007;
temp_data[2910] = 32'h54adaf7d;
temp_data[2911] = 32'h548663e9;
temp_data[2912] = 32'h545af91e;
temp_data[2913] = 32'h542b003f;
temp_data[2914] = 32'h53f5fea0;
temp_data[2915] = 32'h53bb6c2f;
temp_data[2916] = 32'h53843340;
temp_data[2917] = 32'h53522639;
temp_data[2918] = 32'h5324c51e;
temp_data[2919] = 32'h52fb9c41;
temp_data[2920] = 32'h52d642f6;
temp_data[2921] = 32'h52b45a9b;
temp_data[2922] = 32'h52958da4;
temp_data[2923] = 32'h52798ed2;
temp_data[2924] = 32'h52601865;
temp_data[2925] = 32'h5248eb64;
temp_data[2926] = 32'h5233cf07;
temp_data[2927] = 32'h52209019;
temp_data[2928] = 32'h520f0071;
temp_data[2929] = 32'h51fef66f;
temp_data[2930] = 32'h51f04c90;
temp_data[2931] = 32'h51e2e111;
temp_data[2932] = 32'h51d6957d;
temp_data[2933] = 32'h51cb4e62;
temp_data[2934] = 32'h51c0f306;
temp_data[2935] = 32'h51b76d2b;
temp_data[2936] = 32'h51aea8b5;
temp_data[2937] = 32'h51a69392;
temp_data[2938] = 32'h519f1d69;
temp_data[2939] = 32'h51983786;
temp_data[2940] = 32'h5191d4aa;
temp_data[2941] = 32'h518be8d5;
temp_data[2942] = 32'h51866938;
temp_data[2943] = 32'h51814c16;
temp_data[2944] = 32'h517c889c;
temp_data[2945] = 32'h517816db;
temp_data[2946] = 32'h5173ef9a;
temp_data[2947] = 32'h51700c5f;
temp_data[2948] = 32'h516c6745;
temp_data[2949] = 32'h5168faf8;
temp_data[2950] = 32'h5165c2ad;
temp_data[2951] = 32'h5162ba02;
temp_data[2952] = 32'h515fdd05;
temp_data[2953] = 32'h515d2820;
temp_data[2954] = 32'h515a980f;
temp_data[2955] = 32'h515829e1;
temp_data[2956] = 32'h5155dae8;
temp_data[2957] = 32'h5153a8b5;
temp_data[2958] = 32'h5151910c;
temp_data[2959] = 32'h514f91ef;
temp_data[2960] = 32'h514da982;
temp_data[2961] = 32'h514bd61f;
temp_data[2962] = 32'h514a1637;
temp_data[2963] = 32'h5148686a;
temp_data[2964] = 32'h5146cb6c;
temp_data[2965] = 32'h51453e1d;
temp_data[2966] = 32'h5143bf62;
temp_data[2967] = 32'h51424e48;
temp_data[2968] = 32'h5140e9e2;
temp_data[2969] = 32'h513f9164;
temp_data[2970] = 32'h513e440f;
temp_data[2971] = 32'h513d0126;
temp_data[2972] = 32'h513bc811;
temp_data[2973] = 32'h513a982d;
temp_data[2974] = 32'h513970f8;
temp_data[2975] = 32'h513851f0;
temp_data[2976] = 32'h51373a9b;
temp_data[2977] = 32'h51362a8d;
temp_data[2978] = 32'h5135215c;
temp_data[2979] = 32'h51341eac;
temp_data[2980] = 32'h51332225;
temp_data[2981] = 32'h51322b77;
temp_data[2982] = 32'h51313a50;
temp_data[2983] = 32'h51304e6a;
temp_data[2984] = 32'h512f6784;
temp_data[2985] = 32'h512e855e;
temp_data[2986] = 32'h512da7c1;
temp_data[2987] = 32'h512cce74;
temp_data[2988] = 32'h512bf940;
temp_data[2989] = 32'h512b27fa;
temp_data[2990] = 32'h512a5a75;
temp_data[2991] = 32'h51299082;
temp_data[2992] = 32'h5128c9f7;
temp_data[2993] = 32'h512806b3;
temp_data[2994] = 32'h51274691;
temp_data[2995] = 32'h5126896e;
temp_data[2996] = 32'h5125cf29;
temp_data[2997] = 32'h512517a4;
temp_data[2998] = 32'h512462bf;
temp_data[2999] = 32'h5123b060;
temp_data[3000] = 32'h5123006d;
temp_data[3001] = 32'h512252ce;
temp_data[3002] = 32'h5121a769;
temp_data[3003] = 32'h5120fe26;
temp_data[3004] = 32'h512056f3;
temp_data[3005] = 32'h511fb1b8;
temp_data[3006] = 32'h511f0e63;
temp_data[3007] = 32'h511e6cdf;
temp_data[3008] = 32'h511dcd18;
temp_data[3009] = 32'h511d2f01;
temp_data[3010] = 32'h511c9286;
temp_data[3011] = 32'h511bf794;
temp_data[3012] = 32'h511b5e24;
temp_data[3013] = 32'h511ac61e;
temp_data[3014] = 32'h511a2f7b;
temp_data[3015] = 32'h51199a28;
temp_data[3016] = 32'h51190618;
temp_data[3017] = 32'h51187343;
temp_data[3018] = 32'h5117e19c;
temp_data[3019] = 32'h51175111;
temp_data[3020] = 32'h5116c19c;
temp_data[3021] = 32'h51163337;
temp_data[3022] = 32'h5115a5ce;
temp_data[3023] = 32'h5115195d;
temp_data[3024] = 32'h51148dde;
temp_data[3025] = 32'h51140343;
temp_data[3026] = 32'h51137985;
temp_data[3027] = 32'h5112f0a2;
temp_data[3028] = 32'h5112688c;
temp_data[3029] = 32'h5111e143;
temp_data[3030] = 32'h51115abc;
temp_data[3031] = 32'h5110d4f6;
temp_data[3032] = 32'h51104fec;
temp_data[3033] = 32'h510fcb9b;
temp_data[3034] = 32'h510f47fe;
temp_data[3035] = 32'h510ec515;
temp_data[3036] = 32'h510e42e1;
temp_data[3037] = 32'h510dc161;
temp_data[3038] = 32'h510d4096;
temp_data[3039] = 32'h510cc083;
temp_data[3040] = 32'h510c412d;
temp_data[3041] = 32'h510bc298;
temp_data[3042] = 32'h510b44cc;
temp_data[3043] = 32'h510ac7d2;
temp_data[3044] = 32'h510a4bb6;
temp_data[3045] = 32'h5109d081;
temp_data[3046] = 32'h51095647;
temp_data[3047] = 32'h5108dd1a;
temp_data[3048] = 32'h5108650a;
temp_data[3049] = 32'h5107ee35;
temp_data[3050] = 32'h510778b3;
temp_data[3051] = 32'h510704a7;
temp_data[3052] = 32'h51069232;
temp_data[3053] = 32'h5106217d;
temp_data[3054] = 32'h5105b2bc;
temp_data[3055] = 32'h5105461b;
temp_data[3056] = 32'h5104dbdb;
temp_data[3057] = 32'h5104743a;
temp_data[3058] = 32'h51040f88;
temp_data[3059] = 32'h5103ae19;
temp_data[3060] = 32'h51035040;
temp_data[3061] = 32'h5102f673;
temp_data[3062] = 32'h5102a11f;
temp_data[3063] = 32'h510250ca;
temp_data[3064] = 32'h51020608;
temp_data[3065] = 32'h5101c176;
temp_data[3066] = 32'h510183d3;
temp_data[3067] = 32'h51014de4;
temp_data[3068] = 32'h5101208e;
temp_data[3069] = 32'h5100fcd2;
temp_data[3070] = 32'h5100e3c1;
temp_data[3071] = 32'h5100d69d;
temp_data[3072] = 32'h50f6f3a5;
temp_data[3073] = 32'h50f70004;
temp_data[3074] = 32'h50f71783;
temp_data[3075] = 32'h50f738fc;
temp_data[3076] = 32'h50f76352;
temp_data[3077] = 32'h50f7958e;
temp_data[3078] = 32'h50f7ced9;
temp_data[3079] = 32'h50f80e67;
temp_data[3080] = 32'h50f85387;
temp_data[3081] = 32'h50f89d95;
temp_data[3082] = 32'h50f8ec07;
temp_data[3083] = 32'h50f93e5c;
temp_data[3084] = 32'h50f9941d;
temp_data[3085] = 32'h50f9ecea;
temp_data[3086] = 32'h50fa4862;
temp_data[3087] = 32'h50faa633;
temp_data[3088] = 32'h50fb0614;
temp_data[3089] = 32'h50fb67c7;
temp_data[3090] = 32'h50fbcb10;
temp_data[3091] = 32'h50fc2fba;
temp_data[3092] = 32'h50fc9596;
temp_data[3093] = 32'h50fcfc7a;
temp_data[3094] = 32'h50fd6445;
temp_data[3095] = 32'h50fdccd5;
temp_data[3096] = 32'h50fe3611;
temp_data[3097] = 32'h50fe9fd8;
temp_data[3098] = 32'h50ff0a1c;
temp_data[3099] = 32'h50ff74c5;
temp_data[3100] = 32'h50ffdfc2;
temp_data[3101] = 32'h51004b02;
temp_data[3102] = 32'h5100b680;
temp_data[3103] = 32'h51012229;
temp_data[3104] = 32'h51018dfc;
temp_data[3105] = 32'h5101f9e8;
temp_data[3106] = 32'h510265e9;
temp_data[3107] = 32'h5102d1fa;
temp_data[3108] = 32'h51033e18;
temp_data[3109] = 32'h5103aa3b;
temp_data[3110] = 32'h51041666;
temp_data[3111] = 32'h51048295;
temp_data[3112] = 32'h5104eebf;
temp_data[3113] = 32'h51055aee;
temp_data[3114] = 32'h5105c71d;
temp_data[3115] = 32'h5106334c;
temp_data[3116] = 32'h51069f80;
temp_data[3117] = 32'h51070baf;
temp_data[3118] = 32'h510777e6;
temp_data[3119] = 32'h5107e41d;
temp_data[3120] = 32'h51085061;
temp_data[3121] = 32'h5108bca9;
temp_data[3122] = 32'h510928fe;
temp_data[3123] = 32'h51099564;
temp_data[3124] = 32'h510a01d6;
temp_data[3125] = 32'h510a6e5d;
temp_data[3126] = 32'h510adafd;
temp_data[3127] = 32'h510b47b6;
temp_data[3128] = 32'h510bb48d;
temp_data[3129] = 32'h510c2181;
temp_data[3130] = 32'h510c8e9f;
temp_data[3131] = 32'h510cfbe3;
temp_data[3132] = 32'h510d6955;
temp_data[3133] = 32'h510dd6f9;
temp_data[3134] = 32'h510e44d0;
temp_data[3135] = 32'h510eb2dd;
temp_data[3136] = 32'h510f2129;
temp_data[3137] = 32'h510f8fb4;
temp_data[3138] = 32'h510ffe87;
temp_data[3139] = 32'h51106da4;
temp_data[3140] = 32'h5110dd0e;
temp_data[3141] = 32'h51114ccb;
temp_data[3142] = 32'h5111bce0;
temp_data[3143] = 32'h51122d51;
temp_data[3144] = 32'h51129e28;
temp_data[3145] = 32'h51130f5e;
temp_data[3146] = 32'h51138106;
temp_data[3147] = 32'h5113f31b;
temp_data[3148] = 32'h511465a5;
temp_data[3149] = 32'h5114d8ae;
temp_data[3150] = 32'h51154c34;
temp_data[3151] = 32'h5115c040;
temp_data[3152] = 32'h511634db;
temp_data[3153] = 32'h5116aa04;
temp_data[3154] = 32'h51171fc9;
temp_data[3155] = 32'h51179629;
temp_data[3156] = 32'h51180d30;
temp_data[3157] = 32'h511884e0;
temp_data[3158] = 32'h5118fd44;
temp_data[3159] = 32'h5119765c;
temp_data[3160] = 32'h5119f035;
temp_data[3161] = 32'h511a6ad7;
temp_data[3162] = 32'h511ae647;
temp_data[3163] = 32'h511b6289;
temp_data[3164] = 32'h511bdfad;
temp_data[3165] = 32'h511c5db3;
temp_data[3166] = 32'h511cdca9;
temp_data[3167] = 32'h511d5c96;
temp_data[3168] = 32'h511ddd87;
temp_data[3169] = 32'h511e5f81;
temp_data[3170] = 32'h511ee28f;
temp_data[3171] = 32'h511f66ba;
temp_data[3172] = 32'h511fec14;
temp_data[3173] = 32'h5120729f;
temp_data[3174] = 32'h5120fa6a;
temp_data[3175] = 32'h51218384;
temp_data[3176] = 32'h51220dfa;
temp_data[3177] = 32'h512299d9;
temp_data[3178] = 32'h5123272d;
temp_data[3179] = 32'h5123b603;
temp_data[3180] = 32'h5124466f;
temp_data[3181] = 32'h5124d884;
temp_data[3182] = 32'h51256c51;
temp_data[3183] = 32'h512601e2;
temp_data[3184] = 32'h51269952;
temp_data[3185] = 32'h512732b5;
temp_data[3186] = 32'h5127ce1c;
temp_data[3187] = 32'h51286ba0;
temp_data[3188] = 32'h51290b56;
temp_data[3189] = 32'h5129ad5c;
temp_data[3190] = 32'h512a51c6;
temp_data[3191] = 32'h512af8b6;
temp_data[3192] = 32'h512ba240;
temp_data[3193] = 32'h512c4e8b;
temp_data[3194] = 32'h512cfdb1;
temp_data[3195] = 32'h512dafd1;
temp_data[3196] = 32'h512e6517;
temp_data[3197] = 32'h512f1d9f;
temp_data[3198] = 32'h512fd98c;
temp_data[3199] = 32'h5130990b;
temp_data[3200] = 32'h51315c42;
temp_data[3201] = 32'h51322357;
temp_data[3202] = 32'h5132ee74;
temp_data[3203] = 32'h5133bdc7;
temp_data[3204] = 32'h51349175;
temp_data[3205] = 32'h513569ad;
temp_data[3206] = 32'h51364695;
temp_data[3207] = 32'h51372856;
temp_data[3208] = 32'h51380f1f;
temp_data[3209] = 32'h5138fb09;
temp_data[3210] = 32'h5139ec3e;
temp_data[3211] = 32'h513ae2d2;
temp_data[3212] = 32'h513bdee3;
temp_data[3213] = 32'h513ce07a;
temp_data[3214] = 32'h513de79f;
temp_data[3215] = 32'h513ef44d;
temp_data[3216] = 32'h51400670;
temp_data[3217] = 32'h51411deb;
temp_data[3218] = 32'h51423a8a;
temp_data[3219] = 32'h51435c03;
temp_data[3220] = 32'h514481fe;
temp_data[3221] = 32'h5145ac00;
temp_data[3222] = 32'h5146d988;
temp_data[3223] = 32'h514809e1;
temp_data[3224] = 32'h51493c4b;
temp_data[3225] = 32'h514a6feb;
temp_data[3226] = 32'h514ba3c6;
temp_data[3227] = 32'h514cd6d0;
temp_data[3228] = 32'h514e07dd;
temp_data[3229] = 32'h514f3761;
temp_data[3230] = 32'h51506a94;
temp_data[3231] = 32'h5151a049;
temp_data[3232] = 32'h5152d767;
temp_data[3233] = 32'h51540ee9;
temp_data[3234] = 32'h515545ed;
temp_data[3235] = 32'h51567ba6;
temp_data[3236] = 32'h5157af5c;
temp_data[3237] = 32'h5158e083;
temp_data[3238] = 32'h515a0ea2;
temp_data[3239] = 32'h515b3954;
temp_data[3240] = 32'h515c605f;
temp_data[3241] = 32'h515d8390;
temp_data[3242] = 32'h515ea2d3;
temp_data[3243] = 32'h515fbe23;
temp_data[3244] = 32'h5160d584;
temp_data[3245] = 32'h5161e918;
temp_data[3246] = 32'h5162f905;
temp_data[3247] = 32'h51640579;
temp_data[3248] = 32'h51650eb6;
temp_data[3249] = 32'h516614fd;
temp_data[3250] = 32'h516718a4;
temp_data[3251] = 32'h516819fc;
temp_data[3252] = 32'h51691961;
temp_data[3253] = 32'h516a173c;
temp_data[3254] = 32'h516b13f5;
temp_data[3255] = 32'h516c1002;
temp_data[3256] = 32'h516d0bd8;
temp_data[3257] = 32'h516e07ff;
temp_data[3258] = 32'h516f04ff;
temp_data[3259] = 32'h51700368;
temp_data[3260] = 32'h517103de;
temp_data[3261] = 32'h517206ff;
temp_data[3262] = 32'h51730d88;
temp_data[3263] = 32'h5174183b;
temp_data[3264] = 32'h517527e5;
temp_data[3265] = 32'h51763d71;
temp_data[3266] = 32'h517759cd;
temp_data[3267] = 32'h51787e0b;
temp_data[3268] = 32'h5179ab4b;
temp_data[3269] = 32'h517ae2d2;
temp_data[3270] = 32'h517c25f6;
temp_data[3271] = 32'h517d7642;
temp_data[3272] = 32'h517ed552;
temp_data[3273] = 32'h518044fe;
temp_data[3274] = 32'h5181c73b;
temp_data[3275] = 32'h51835e4a;
temp_data[3276] = 32'h51850c91;
temp_data[3277] = 32'h5186d4c3;
temp_data[3278] = 32'h5188b9d8;
temp_data[3279] = 32'h518abf23;
temp_data[3280] = 32'h518ce847;
temp_data[3281] = 32'h518f3950;
temp_data[3282] = 32'h5191b6bb;
temp_data[3283] = 32'h51946584;
temp_data[3284] = 32'h51974b38;
temp_data[3285] = 32'h519a6df0;
temp_data[3286] = 32'h519dd484;
temp_data[3287] = 32'h51a18683;
temp_data[3288] = 32'h51a58c54;
temp_data[3289] = 32'h51a9ef46;
temp_data[3290] = 32'h51aeb9b6;
temp_data[3291] = 32'h51b3f71f;
temp_data[3292] = 32'h51b9b439;
temp_data[3293] = 32'h51bfff1e;
temp_data[3294] = 32'h51c6e771;
temp_data[3295] = 32'h51ce7e74;
temp_data[3296] = 32'h51d6d745;
temp_data[3297] = 32'h51e00707;
temp_data[3298] = 32'h51ea2503;
temp_data[3299] = 32'h51f54b12;
temp_data[3300] = 32'h51ffbe98;
temp_data[3301] = 32'h52092489;
temp_data[3302] = 32'h521194af;
temp_data[3303] = 32'h5219245b;
temp_data[3304] = 32'h521fe675;
temp_data[3305] = 32'h5225ebc8;
temp_data[3306] = 32'h522b4313;
temp_data[3307] = 32'h522ff940;
temp_data[3308] = 32'h52341976;
temp_data[3309] = 32'h5237ad36;
temp_data[3310] = 32'h523abc84;
temp_data[3311] = 32'h523d4de4;
temp_data[3312] = 32'h523f6680;
temp_data[3313] = 32'h52410a28;
temp_data[3314] = 32'h52423b75;
temp_data[3315] = 32'h5242fbb5;
temp_data[3316] = 32'h52434afd;
temp_data[3317] = 32'h52432831;
temp_data[3318] = 32'h52429100;
temp_data[3319] = 32'h524181d8;
temp_data[3320] = 32'h523ff5e0;
temp_data[3321] = 32'h523de6ff;
temp_data[3322] = 32'h523b4db6;
temp_data[3323] = 32'h52382110;
temp_data[3324] = 32'h523456ac;
temp_data[3325] = 32'h522fe271;
temp_data[3326] = 32'h522ab69a;
temp_data[3327] = 32'h5224c383;
temp_data[3328] = 32'h521df762;
temp_data[3329] = 32'h521813db;
temp_data[3330] = 32'h5213073e;
temp_data[3331] = 32'h520ec212;
temp_data[3332] = 32'h520b36d6;
temp_data[3333] = 32'h520859e6;
temp_data[3334] = 32'h5206214b;
temp_data[3335] = 32'h520484b6;
temp_data[3336] = 32'h52037d56;
temp_data[3337] = 32'h520305e6;
temp_data[3338] = 32'h52031a7e;
temp_data[3339] = 32'h5203b8aa;
temp_data[3340] = 32'h5204df4c;
temp_data[3341] = 32'h52068eb0;
temp_data[3342] = 32'h5208c87e;
temp_data[3343] = 32'h520b8fc9;
temp_data[3344] = 32'h520ee910;
temp_data[3345] = 32'h5212da62;
temp_data[3346] = 32'h52176b51;
temp_data[3347] = 32'h521ca527;
temp_data[3348] = 32'h522292ea;
temp_data[3349] = 32'h52294189;
temp_data[3350] = 32'h5230c001;
temp_data[3351] = 32'h52391f82;
temp_data[3352] = 32'h524273a3;
temp_data[3353] = 32'h524cd2a2;
temp_data[3354] = 32'h5258559b;
temp_data[3355] = 32'h526518ce;
temp_data[3356] = 32'h52733bf7;
temp_data[3357] = 32'h5282e2a4;
temp_data[3358] = 32'h52943498;
temp_data[3359] = 32'h52a75e31;
temp_data[3360] = 32'h52bc90fb;
temp_data[3361] = 32'h52d40410;
temp_data[3362] = 32'h52edf4cf;
temp_data[3363] = 32'h530aa769;
temp_data[3364] = 32'h532a678c;
temp_data[3365] = 32'h534d8933;
temp_data[3366] = 32'h5374696a;
temp_data[3367] = 32'h539f6f33;
temp_data[3368] = 32'h53cf0c84;
temp_data[3369] = 32'h5403bf94;
temp_data[3370] = 32'h54398030;
temp_data[3371] = 32'h5469fef4;
temp_data[3372] = 32'h5495bcba;
temp_data[3373] = 32'h54bd2dba;
temp_data[3374] = 32'h54e0bafe;
temp_data[3375] = 32'h5500c365;
temp_data[3376] = 32'h551d9c88;
temp_data[3377] = 32'h5537938a;
temp_data[3378] = 32'h554eede5;
temp_data[3379] = 32'h5563ea14;
temp_data[3380] = 32'h5576c02b;
temp_data[3381] = 32'h5587a287;
temp_data[3382] = 32'h5596be40;
temp_data[3383] = 32'h55a43bb0;
temp_data[3384] = 32'h55b03ed1;
temp_data[3385] = 32'h55bae7c0;
temp_data[3386] = 32'h55c452fc;
temp_data[3387] = 32'h55cc99bf;
temp_data[3388] = 32'h55d3d252;
temp_data[3389] = 32'h55da1038;
temp_data[3390] = 32'h55df647c;
temp_data[3391] = 32'h55e3ddd3;
temp_data[3392] = 32'h55e788c2;
temp_data[3393] = 32'h55ea6fdf;
temp_data[3394] = 32'h55ec9bc7;
temp_data[3395] = 32'h55ee135e;
temp_data[3396] = 32'h55eedbc6;
temp_data[3397] = 32'h55eef883;
temp_data[3398] = 32'h55ee6b72;
temp_data[3399] = 32'h55ed34e3;
temp_data[3400] = 32'h55eb5382;
temp_data[3401] = 32'h55e8c476;
temp_data[3402] = 32'h55e58334;
temp_data[3403] = 32'h55e18987;
temp_data[3404] = 32'h55dccf7d;
temp_data[3405] = 32'h55d74b49;
temp_data[3406] = 32'h55d0f135;
temp_data[3407] = 32'h55c9b368;
temp_data[3408] = 32'h55c181dc;
temp_data[3409] = 32'h55b84a1b;
temp_data[3410] = 32'h55adf712;
temp_data[3411] = 32'h55a270d6;
temp_data[3412] = 32'h55959c52;
temp_data[3413] = 32'h55875b18;
temp_data[3414] = 32'h55778ae7;
temp_data[3415] = 32'h55660568;
temp_data[3416] = 32'h55529fb6;
temp_data[3417] = 32'h553d29e1;
temp_data[3418] = 32'h55256e7a;
temp_data[3419] = 32'h550b31fd;
temp_data[3420] = 32'h54ee3227;
temp_data[3421] = 32'h54ce255b;
temp_data[3422] = 32'h54aab9e5;
temp_data[3423] = 32'h5483951c;
temp_data[3424] = 32'h5458528b;
temp_data[3425] = 32'h54288302;
temp_data[3426] = 32'h53f3ab71;
temp_data[3427] = 32'h53b9435f;
temp_data[3428] = 32'h538234b9;
temp_data[3429] = 32'h53505172;
temp_data[3430] = 32'h5323192f;
temp_data[3431] = 32'h52fa17e7;
temp_data[3432] = 32'h52d4e4a4;
temp_data[3433] = 32'h52b32086;
temp_data[3434] = 32'h529475cd;
temp_data[3435] = 32'h52789720;
temp_data[3436] = 32'h525f3ea7;
temp_data[3437] = 32'h52482d66;
temp_data[3438] = 32'h52332a9d;
temp_data[3439] = 32'h52200321;
temp_data[3440] = 32'h520e88db;
temp_data[3441] = 32'h51fe924b;
temp_data[3442] = 32'h51effa09;
temp_data[3443] = 32'h51e29e67;
temp_data[3444] = 32'h51d66117;
temp_data[3445] = 32'h51cb26c8;
temp_data[3446] = 32'h51c0d6e0;
temp_data[3447] = 32'h51b75b36;
temp_data[3448] = 32'h51ae9fcf;
temp_data[3449] = 32'h51a692b0;
temp_data[3450] = 32'h519f23a3;
temp_data[3451] = 32'h51984403;
temp_data[3452] = 32'h5191e6a3;
temp_data[3453] = 32'h518bffa0;
temp_data[3454] = 32'h5186843c;
temp_data[3455] = 32'h51816ac2;
temp_data[3456] = 32'h517caa7a;
temp_data[3457] = 32'h51783b71;
temp_data[3458] = 32'h5174168b;
temp_data[3459] = 32'h51703550;
temp_data[3460] = 32'h516c91e6;
temp_data[3461] = 32'h51692707;
temp_data[3462] = 32'h5165efe5;
temp_data[3463] = 32'h5162e82d;
temp_data[3464] = 32'h51600bf6;
temp_data[3465] = 32'h515d57a3;
temp_data[3466] = 32'h515ac804;
temp_data[3467] = 32'h51585a25;
temp_data[3468] = 32'h51560b5f;
temp_data[3469] = 32'h5153d940;
temp_data[3470] = 32'h5151c194;
temp_data[3471] = 32'h514fc261;
temp_data[3472] = 32'h514dd9cb;
temp_data[3473] = 32'h514c0629;
temp_data[3474] = 32'h514a45fa;
temp_data[3475] = 32'h514897d9;
temp_data[3476] = 32'h5146fa7f;
temp_data[3477] = 32'h51456cc2;
temp_data[3478] = 32'h5143ed9a;
temp_data[3479] = 32'h51427c03;
temp_data[3480] = 32'h51411722;
temp_data[3481] = 32'h513fbe23;
temp_data[3482] = 32'h513e703f;
temp_data[3483] = 32'h513d2ccf;
temp_data[3484] = 32'h513bf328;
temp_data[3485] = 32'h513ac2b5;
temp_data[3486] = 32'h51399aed;
temp_data[3487] = 32'h51387b4e;
temp_data[3488] = 32'h5137635e;
temp_data[3489] = 32'h513652b9;
temp_data[3490] = 32'h513548ed;
temp_data[3491] = 32'h513445a6;
temp_data[3492] = 32'h51334884;
temp_data[3493] = 32'h51325137;
temp_data[3494] = 32'h51315f78;
temp_data[3495] = 32'h513072f7;
temp_data[3496] = 32'h512f8b76;
temp_data[3497] = 32'h512ea8b9;
temp_data[3498] = 32'h512dca82;
temp_data[3499] = 32'h512cf099;
temp_data[3500] = 32'h512c1ad2;
temp_data[3501] = 32'h512b48f5;
temp_data[3502] = 32'h512a7ad5;
temp_data[3503] = 32'h5129b04f;
temp_data[3504] = 32'h5128e932;
temp_data[3505] = 32'h51282557;
temp_data[3506] = 32'h512764a1;
temp_data[3507] = 32'h5126a6ec;
temp_data[3508] = 32'h5125ec14;
temp_data[3509] = 32'h51253401;
temp_data[3510] = 32'h51247e8d;
temp_data[3511] = 32'h5123cb9f;
temp_data[3512] = 32'h51231b1e;
temp_data[3513] = 32'h51226cf4;
temp_data[3514] = 32'h5121c101;
temp_data[3515] = 32'h51211737;
temp_data[3516] = 32'h51206f7a;
temp_data[3517] = 32'h511fc9b4;
temp_data[3518] = 32'h511f25d9;
temp_data[3519] = 32'h511e83cb;
temp_data[3520] = 32'h511de382;
temp_data[3521] = 32'h511d44e5;
temp_data[3522] = 32'h511ca7e3;
temp_data[3523] = 32'h511c0c74;
temp_data[3524] = 32'h511b727e;
temp_data[3525] = 32'h511ad9f9;
temp_data[3526] = 32'h511a42d5;
temp_data[3527] = 32'h5119ad00;
temp_data[3528] = 32'h51191876;
temp_data[3529] = 32'h51188523;
temp_data[3530] = 32'h5117f2fa;
temp_data[3531] = 32'h511761f6;
temp_data[3532] = 32'h5116d207;
temp_data[3533] = 32'h51164324;
temp_data[3534] = 32'h5115b542;
temp_data[3535] = 32'h5115285b;
temp_data[3536] = 32'h51149c63;
temp_data[3537] = 32'h51141151;
temp_data[3538] = 32'h5113871e;
temp_data[3539] = 32'h5112fdc1;
temp_data[3540] = 32'h5112753a;
temp_data[3541] = 32'h5111ed78;
temp_data[3542] = 32'h51116680;
temp_data[3543] = 32'h5110e048;
temp_data[3544] = 32'h51105acd;
temp_data[3545] = 32'h510fd60a;
temp_data[3546] = 32'h510f51fc;
temp_data[3547] = 32'h510ecea7;
temp_data[3548] = 32'h510e4c06;
temp_data[3549] = 32'h510dca19;
temp_data[3550] = 32'h510d48e0;
temp_data[3551] = 32'h510cc865;
temp_data[3552] = 32'h510c48a1;
temp_data[3553] = 32'h510bc9a3;
temp_data[3554] = 32'h510b4b6f;
temp_data[3555] = 32'h510ace10;
temp_data[3556] = 32'h510a518b;
temp_data[3557] = 32'h5109d5f5;
temp_data[3558] = 32'h51095b57;
temp_data[3559] = 32'h5108e1c6;
temp_data[3560] = 32'h51086955;
temp_data[3561] = 32'h5107f224;
temp_data[3562] = 32'h51077c42;
temp_data[3563] = 32'h510707d9;
temp_data[3564] = 32'h5106950c;
temp_data[3565] = 32'h510623ff;
temp_data[3566] = 32'h5105b4e5;
temp_data[3567] = 32'h510547f5;
temp_data[3568] = 32'h5104dd61;
temp_data[3569] = 32'h51047575;
temp_data[3570] = 32'h51041077;
temp_data[3571] = 32'h5103aebc;
temp_data[3572] = 32'h510350a0;
temp_data[3573] = 32'h5102f690;
temp_data[3574] = 32'h5102a101;
temp_data[3575] = 32'h51025072;
temp_data[3576] = 32'h51020579;
temp_data[3577] = 32'h5101c0be;
temp_data[3578] = 32'h510182ed;
temp_data[3579] = 32'h51014cdb;
temp_data[3580] = 32'h51011f6d;
temp_data[3581] = 32'h5100fb98;
temp_data[3582] = 32'h5100e27a;
temp_data[3583] = 32'h5100d54e;
temp_data[3584] = 32'h50f6e8e6;
temp_data[3585] = 32'h50f6f549;
temp_data[3586] = 32'h50f70cd4;
temp_data[3587] = 32'h50f72e5e;
temp_data[3588] = 32'h50f758c9;
temp_data[3589] = 32'h50f78b26;
temp_data[3590] = 32'h50f7c48f;
temp_data[3591] = 32'h50f80443;
temp_data[3592] = 32'h50f84990;
temp_data[3593] = 32'h50f893d1;
temp_data[3594] = 32'h50f8e27a;
temp_data[3595] = 32'h50f93505;
temp_data[3596] = 32'h50f98b05;
temp_data[3597] = 32'h50f9e411;
temp_data[3598] = 32'h50fa3fcd;
temp_data[3599] = 32'h50fa9de5;
temp_data[3600] = 32'h50fafe11;
temp_data[3601] = 32'h50fb600f;
temp_data[3602] = 32'h50fbc3a8;
temp_data[3603] = 32'h50fc28a2;
temp_data[3604] = 32'h50fc8ed2;
temp_data[3605] = 32'h50fcf60a;
temp_data[3606] = 32'h50fd5e2d;
temp_data[3607] = 32'h50fdc715;
temp_data[3608] = 32'h50fe30a9;
temp_data[3609] = 32'h50fe9acc;
temp_data[3610] = 32'h50ff056c;
temp_data[3611] = 32'h50ff7072;
temp_data[3612] = 32'h50ffdbcf;
temp_data[3613] = 32'h51004773;
temp_data[3614] = 32'h5100b34e;
temp_data[3615] = 32'h51011f5c;
temp_data[3616] = 32'h51018b8f;
temp_data[3617] = 32'h5101f7e0;
temp_data[3618] = 32'h51026445;
temp_data[3619] = 32'h5102d0bb;
temp_data[3620] = 32'h51033d3e;
temp_data[3621] = 32'h5103a9ce;
temp_data[3622] = 32'h5104165d;
temp_data[3623] = 32'h510482f5;
temp_data[3624] = 32'h5104ef8d;
temp_data[3625] = 32'h51055c25;
temp_data[3626] = 32'h5105c8bd;
temp_data[3627] = 32'h51063559;
temp_data[3628] = 32'h5106a1f5;
temp_data[3629] = 32'h51070e91;
temp_data[3630] = 32'h51077b35;
temp_data[3631] = 32'h5107e7da;
temp_data[3632] = 32'h5108548b;
temp_data[3633] = 32'h5108c140;
temp_data[3634] = 32'h51092e06;
temp_data[3635] = 32'h51099ad8;
temp_data[3636] = 32'h510a07bc;
temp_data[3637] = 32'h510a74b4;
temp_data[3638] = 32'h510ae1c6;
temp_data[3639] = 32'h510b4ef0;
temp_data[3640] = 32'h510bbc38;
temp_data[3641] = 32'h510c29a6;
temp_data[3642] = 32'h510c9735;
temp_data[3643] = 32'h510d04ee;
temp_data[3644] = 32'h510d72d6;
temp_data[3645] = 32'h510de0eb;
temp_data[3646] = 32'h510e4f3c;
temp_data[3647] = 32'h510ebdbe;
temp_data[3648] = 32'h510f2c84;
temp_data[3649] = 32'h510f9b89;
temp_data[3650] = 32'h51100ad4;
temp_data[3651] = 32'h51107a6c;
temp_data[3652] = 32'h5110ea4f;
temp_data[3653] = 32'h51115a8a;
temp_data[3654] = 32'h5111cb1d;
temp_data[3655] = 32'h51123c0c;
temp_data[3656] = 32'h5112ad5c;
temp_data[3657] = 32'h51131f15;
temp_data[3658] = 32'h5113913a;
temp_data[3659] = 32'h511403d1;
temp_data[3660] = 32'h511476de;
temp_data[3661] = 32'h5114ea68;
temp_data[3662] = 32'h51155e74;
temp_data[3663] = 32'h5115d307;
temp_data[3664] = 32'h51164828;
temp_data[3665] = 32'h5116bddc;
temp_data[3666] = 32'h51173426;
temp_data[3667] = 32'h5117ab11;
temp_data[3668] = 32'h511822a3;
temp_data[3669] = 32'h51189ae1;
temp_data[3670] = 32'h511913d3;
temp_data[3671] = 32'h51198d7e;
temp_data[3672] = 32'h511a07ea;
temp_data[3673] = 32'h511a831b;
temp_data[3674] = 32'h511aff22;
temp_data[3675] = 32'h511b7bfa;
temp_data[3676] = 32'h511bf9b5;
temp_data[3677] = 32'h511c785b;
temp_data[3678] = 32'h511cf7f0;
temp_data[3679] = 32'h511d787d;
temp_data[3680] = 32'h511dfa0d;
temp_data[3681] = 32'h511e7caf;
temp_data[3682] = 32'h511f0065;
temp_data[3683] = 32'h511f853c;
temp_data[3684] = 32'h51200b41;
temp_data[3685] = 32'h5120927d;
temp_data[3686] = 32'h51211b00;
temp_data[3687] = 32'h5121a4d3;
temp_data[3688] = 32'h51223006;
temp_data[3689] = 32'h5122bca5;
temp_data[3690] = 32'h51234abe;
temp_data[3691] = 32'h5123da62;
temp_data[3692] = 32'h51246ba0;
temp_data[3693] = 32'h5124fe8b;
temp_data[3694] = 32'h51259336;
temp_data[3695] = 32'h512629ae;
temp_data[3696] = 32'h5126c209;
temp_data[3697] = 32'h51275c5f;
temp_data[3698] = 32'h5127f8c6;
temp_data[3699] = 32'h51289753;
temp_data[3700] = 32'h5129381d;
temp_data[3701] = 32'h5129db44;
temp_data[3702] = 32'h512a80dc;
temp_data[3703] = 32'h512b2907;
temp_data[3704] = 32'h512bd3e1;
temp_data[3705] = 32'h512c8188;
temp_data[3706] = 32'h512d3223;
temp_data[3707] = 32'h512de5cd;
temp_data[3708] = 32'h512e9cb2;
temp_data[3709] = 32'h512f56f3;
temp_data[3710] = 32'h513014be;
temp_data[3711] = 32'h5130d639;
temp_data[3712] = 32'h51319b8d;
temp_data[3713] = 32'h513264e9;
temp_data[3714] = 32'h5133327b;
temp_data[3715] = 32'h51340471;
temp_data[3716] = 32'h5134daf9;
temp_data[3717] = 32'h5135b64a;
temp_data[3718] = 32'h5136968d;
temp_data[3719] = 32'h51377bf6;
temp_data[3720] = 32'h513866ae;
temp_data[3721] = 32'h513956e7;
temp_data[3722] = 32'h513a4ccb;
temp_data[3723] = 32'h513b4877;
temp_data[3724] = 32'h513c4a12;
temp_data[3725] = 32'h513d51b1;
temp_data[3726] = 32'h513e5f67;
temp_data[3727] = 32'h513f7332;
temp_data[3728] = 32'h51408d0d;
temp_data[3729] = 32'h5141acde;
temp_data[3730] = 32'h5142d27c;
temp_data[3731] = 32'h5143fda0;
temp_data[3732] = 32'h51452df1;
temp_data[3733] = 32'h514662fe;
temp_data[3734] = 32'h51479c34;
temp_data[3735] = 32'h5148d8dc;
temp_data[3736] = 32'h514a182b;
temp_data[3737] = 32'h514b5929;
temp_data[3738] = 32'h514c9acc;
temp_data[3739] = 32'h514ddbe4;
temp_data[3740] = 32'h514f1b33;
temp_data[3741] = 32'h515058fb;
temp_data[3742] = 32'h51519a5b;
temp_data[3743] = 32'h5152de01;
temp_data[3744] = 32'h515422bc;
temp_data[3745] = 32'h51556766;
temp_data[3746] = 32'h5156ab0d;
temp_data[3747] = 32'h5157ecc8;
temp_data[3748] = 32'h51592bdc;
temp_data[3749] = 32'h515a67b6;
temp_data[3750] = 32'h515b9fcf;
temp_data[3751] = 32'h515cd3d4;
temp_data[3752] = 32'h515e0382;
temp_data[3753] = 32'h515f2eb2;
temp_data[3754] = 32'h51605550;
temp_data[3755] = 32'h51617760;
temp_data[3756] = 32'h516294f7;
temp_data[3757] = 32'h5163ae36;
temp_data[3758] = 32'h5164c350;
temp_data[3759] = 32'h5165d480;
temp_data[3760] = 32'h5166e211;
temp_data[3761] = 32'h5167ec46;
temp_data[3762] = 32'h5168f380;
temp_data[3763] = 32'h5169f816;
temp_data[3764] = 32'h516afa6e;
temp_data[3765] = 32'h516bfaf4;
temp_data[3766] = 32'h516cfa16;
temp_data[3767] = 32'h516df851;
temp_data[3768] = 32'h516ef61b;
temp_data[3769] = 32'h516ff402;
temp_data[3770] = 32'h5170f288;
temp_data[3771] = 32'h5171f252;
temp_data[3772] = 32'h5172f3f1;
temp_data[3773] = 32'h5173f81a;
temp_data[3774] = 32'h5174ff7a;
temp_data[3775] = 32'h51760add;
temp_data[3776] = 32'h51771b0d;
temp_data[3777] = 32'h517830f0;
temp_data[3778] = 32'h51794d7f;
temp_data[3779] = 32'h517a71c1;
temp_data[3780] = 32'h517b9edc;
temp_data[3781] = 32'h517cd60f;
temp_data[3782] = 32'h517e18b1;
temp_data[3783] = 32'h517f6840;
temp_data[3784] = 32'h5180c661;
temp_data[3785] = 32'h518234df;
temp_data[3786] = 32'h5183b5b7;
temp_data[3787] = 32'h51854b1b;
temp_data[3788] = 32'h5186f76a;
temp_data[3789] = 32'h5188bd5a;
temp_data[3790] = 32'h518a9fdc;
temp_data[3791] = 32'h518ca234;
temp_data[3792] = 32'h518ec800;
temp_data[3793] = 32'h51911548;
temp_data[3794] = 32'h51938e7e;
temp_data[3795] = 32'h5196389b;
temp_data[3796] = 32'h5199191a;
temp_data[3797] = 32'h519c3615;
temp_data[3798] = 32'h519f9657;
temp_data[3799] = 32'h51a34168;
temp_data[3800] = 32'h51a73fab;
temp_data[3801] = 32'h51ab9a70;
temp_data[3802] = 32'h51b05c07;
temp_data[3803] = 32'h51b58ff3;
temp_data[3804] = 32'h51bb42f6;
temp_data[3805] = 32'h51c1832c;
temp_data[3806] = 32'h51c86042;
temp_data[3807] = 32'h51cfeb9e;
temp_data[3808] = 32'h51d83869;
temp_data[3809] = 32'h51e15be6;
temp_data[3810] = 32'h51eb6d83;
temp_data[3811] = 32'h51f68733;
temp_data[3812] = 32'h5200ee8d;
temp_data[3813] = 32'h520a489d;
temp_data[3814] = 32'h5212ad58;
temp_data[3815] = 32'h521a3223;
temp_data[3816] = 32'h5220ea0c;
temp_data[3817] = 32'h5226e5e6;
temp_data[3818] = 32'h522c348f;
temp_data[3819] = 32'h5230e2ef;
temp_data[3820] = 32'h5234fc37;
temp_data[3821] = 32'h523889f0;
temp_data[3822] = 32'h523b9410;
temp_data[3823] = 32'h523e2121;
temp_data[3824] = 32'h5240363b;
temp_data[3825] = 32'h5241d734;
temp_data[3826] = 32'h5243068e;
temp_data[3827] = 32'h5243c58b;
temp_data[3828] = 32'h52441440;
temp_data[3829] = 32'h5243f17c;
temp_data[3830] = 32'h52435ade;
temp_data[3831] = 32'h52424ccb;
temp_data[3832] = 32'h5240c25d;
temp_data[3833] = 32'h523eb56c;
temp_data[3834] = 32'h523c1e69;
temp_data[3835] = 32'h5238f45a;
temp_data[3836] = 32'h52352cc3;
temp_data[3837] = 32'h5230bb88;
temp_data[3838] = 32'h522b92d5;
temp_data[3839] = 32'h5225a2f0;
temp_data[3840] = 32'h521eda0a;
temp_data[3841] = 32'h5218f9ad;
temp_data[3842] = 32'h5213f028;
temp_data[3843] = 32'h520fadef;
temp_data[3844] = 32'h520c2570;
temp_data[3845] = 32'h52094af9;
temp_data[3846] = 32'h52071487;
temp_data[3847] = 32'h520579b7;
temp_data[3848] = 32'h520473b0;
temp_data[3849] = 32'h5203fd11;
temp_data[3850] = 32'h520411ed;
temp_data[3851] = 32'h5204afb8;
temp_data[3852] = 32'h5205d549;
temp_data[3853] = 32'h520782cf;
temp_data[3854] = 32'h5209b9e5;
temp_data[3855] = 32'h520c7d80;
temp_data[3856] = 32'h520fd21c;
temp_data[3857] = 32'h5213bd98;
temp_data[3858] = 32'h5218477c;
temp_data[3859] = 32'h521d78f2;
temp_data[3860] = 32'h52235ce2;
temp_data[3861] = 32'h522a0022;
temp_data[3862] = 32'h52317182;
temp_data[3863] = 32'h5239c216;
temp_data[3864] = 32'h52430557;
temp_data[3865] = 32'h524d5155;
temp_data[3866] = 32'h5258bf05;
temp_data[3867] = 32'h52656a8c;
temp_data[3868] = 32'h52737375;
temp_data[3869] = 32'h5282fd33;
temp_data[3870] = 32'h52942f6a;
temp_data[3871] = 32'h52a73665;
temp_data[3872] = 32'h52bc439a;
temp_data[3873] = 32'h52d38e22;
temp_data[3874] = 32'h52ed5365;
temp_data[3875] = 32'h5309d7aa;
temp_data[3876] = 32'h532966d3;
temp_data[3877] = 32'h534c5515;
temp_data[3878] = 32'h5372ffd6;
temp_data[3879] = 32'h539dce7d;
temp_data[3880] = 32'h53cd3376;
temp_data[3881] = 32'h5401ad86;
temp_data[3882] = 32'h54373505;
temp_data[3883] = 32'h54677b20;
temp_data[3884] = 32'h54930132;
temp_data[3885] = 32'h54ba3bf7;
temp_data[3886] = 32'h54dd94e2;
temp_data[3887] = 32'h54fd6b2b;
temp_data[3888] = 32'h551a14ad;
temp_data[3889] = 32'h5533dec6;
temp_data[3890] = 32'h554b0f02;
temp_data[3891] = 32'h555fe3eb;
temp_data[3892] = 32'h5572959a;
temp_data[3893] = 32'h55835660;
temp_data[3894] = 32'h55925337;
temp_data[3895] = 32'h559fb463;
temp_data[3896] = 32'h55ab9dc3;
temp_data[3897] = 32'h55b62f4d;
temp_data[3898] = 32'h55bf8559;
temp_data[3899] = 32'h55c7b90a;
temp_data[3900] = 32'h55cee07a;
temp_data[3901] = 32'h55d50f17;
temp_data[3902] = 32'h55da55c5;
temp_data[3903] = 32'h55dec322;
temp_data[3904] = 32'h55e2639d;
temp_data[3905] = 32'h55e541af;
temp_data[3906] = 32'h55e765ed;
temp_data[3907] = 32'h55e8d723;
temp_data[3908] = 32'h55e99a70;
temp_data[3909] = 32'h55e9b342;
temp_data[3910] = 32'h55e92379;
temp_data[3911] = 32'h55e7eb5b;
temp_data[3912] = 32'h55e609a6;
temp_data[3913] = 32'h55e37b70;
temp_data[3914] = 32'h55e03c43;
temp_data[3915] = 32'h55dc45ed;
temp_data[3916] = 32'h55d79093;
temp_data[3917] = 32'h55d2126f;
temp_data[3918] = 32'h55cbbfe4;
temp_data[3919] = 32'h55c48b33;
temp_data[3920] = 32'h55bc646f;
temp_data[3921] = 32'h55b3393b;
temp_data[3922] = 32'h55a8f4a5;
temp_data[3923] = 32'h559d7ee5;
temp_data[3924] = 32'h5590bd0e;
temp_data[3925] = 32'h558290cd;
temp_data[3926] = 32'h5572d806;
temp_data[3927] = 32'h55616c87;
temp_data[3928] = 32'h554e2379;
temp_data[3929] = 32'h5538cd10;
temp_data[3930] = 32'h552133df;
temp_data[3931] = 32'h55071c65;
temp_data[3932] = 32'h54ea4456;
temp_data[3933] = 32'h54ca61f6;
temp_data[3934] = 32'h54a72360;
temp_data[3935] = 32'h54802d9d;
temp_data[3936] = 32'h54551beb;
temp_data[3937] = 32'h54257eaa;
temp_data[3938] = 32'h53f0da51;
temp_data[3939] = 32'h53b6a5db;
temp_data[3940] = 32'h537fcaac;
temp_data[3941] = 32'h534e1a37;
temp_data[3942] = 32'h53211398;
temp_data[3943] = 32'h52f8425f;
temp_data[3944] = 32'h52d33d29;
temp_data[3945] = 32'h52b1a4cf;
temp_data[3946] = 32'h52932360;
temp_data[3947] = 32'h52776b55;
temp_data[3948] = 32'h525e36c6;
temp_data[3949] = 32'h524746bb;
temp_data[3950] = 32'h5232627c;
temp_data[3951] = 32'h521f56eb;
temp_data[3952] = 32'h520df616;
temp_data[3953] = 32'h51fe1694;
temp_data[3954] = 32'h51ef932d;
temp_data[3955] = 32'h51e24a56;
temp_data[3956] = 32'h51d61de2;
temp_data[3957] = 32'h51caf2b2;
temp_data[3958] = 32'h51c0b047;
temp_data[3959] = 32'h51b7409e;
temp_data[3960] = 32'h51ae8feb;
temp_data[3961] = 32'h51a68c43;
temp_data[3962] = 32'h519f2596;
temp_data[3963] = 32'h51984d5e;
temp_data[3964] = 32'h5191f67f;
temp_data[3965] = 32'h518c152f;
temp_data[3966] = 32'h51869ec7;
temp_data[3967] = 32'h518189a9;
temp_data[3968] = 32'h517ccd25;
temp_data[3969] = 32'h51786163;
temp_data[3970] = 32'h51743f4f;
temp_data[3971] = 32'h5170607c;
temp_data[3972] = 32'h516cbf1f;
temp_data[3973] = 32'h516955f8;
temp_data[3974] = 32'h51662047;
temp_data[3975] = 32'h516319c1;
temp_data[3976] = 32'h51603e79;
temp_data[3977] = 32'h515d8af0;
temp_data[3978] = 32'h515afbe3;
temp_data[3979] = 32'h51588e71;
temp_data[3980] = 32'h51563ff2;
temp_data[3981] = 32'h51540dfe;
temp_data[3982] = 32'h5151f666;
temp_data[3983] = 32'h514ff723;
temp_data[3984] = 32'h514e0e6f;
temp_data[3985] = 32'h514c3a9b;
temp_data[3986] = 32'h514a7a29;
temp_data[3987] = 32'h5148cbb4;
temp_data[3988] = 32'h51472dfd;
temp_data[3989] = 32'h51459fd8;
temp_data[3990] = 32'h5144203a;
temp_data[3991] = 32'h5142ae29;
temp_data[3992] = 32'h514148c3;
temp_data[3993] = 32'h513fef39;
temp_data[3994] = 32'h513ea0c7;
temp_data[3995] = 32'h513d5cc0;
temp_data[3996] = 32'h513c2281;
temp_data[3997] = 32'h513af16f;
temp_data[3998] = 32'h5139c908;
temp_data[3999] = 32'h5138a8ca;
temp_data[4000] = 32'h5137903a;
temp_data[4001] = 32'h51367eed;
temp_data[4002] = 32'h5135747e;
temp_data[4003] = 32'h5134708f;
temp_data[4004] = 32'h513372c5;
temp_data[4005] = 32'h51327ad1;
temp_data[4006] = 32'h51318866;
temp_data[4007] = 32'h51309b41;
temp_data[4008] = 32'h512fb318;
temp_data[4009] = 32'h512ecfb3;
temp_data[4010] = 32'h512df0d4;
temp_data[4011] = 32'h512d1644;
temp_data[4012] = 32'h512c3fd5;
temp_data[4013] = 32'h512b6d55;
temp_data[4014] = 32'h512a9e90;
temp_data[4015] = 32'h5129d363;
temp_data[4016] = 32'h51290ba2;
temp_data[4017] = 32'h51284728;
temp_data[4018] = 32'h512785d3;
temp_data[4019] = 32'h5126c77a;
temp_data[4020] = 32'h51260c02;
temp_data[4021] = 32'h51255350;
temp_data[4022] = 32'h51249d3d;
temp_data[4023] = 32'h5123e9b4;
temp_data[4024] = 32'h5123389b;
temp_data[4025] = 32'h512289d2;
temp_data[4026] = 32'h5121dd48;
temp_data[4027] = 32'h512132e4;
temp_data[4028] = 32'h51208a8f;
temp_data[4029] = 32'h511fe436;
temp_data[4030] = 32'h511f3fc4;
temp_data[4031] = 32'h511e9d24;
temp_data[4032] = 32'h511dfc44;
temp_data[4033] = 32'h511d5d18;
temp_data[4034] = 32'h511cbf87;
temp_data[4035] = 32'h511c2381;
temp_data[4036] = 32'h511b8901;
temp_data[4037] = 32'h511aefed;
temp_data[4038] = 32'h511a583a;
temp_data[4039] = 32'h5119c1db;
temp_data[4040] = 32'h51192cc3;
temp_data[4041] = 32'h511898e5;
temp_data[4042] = 32'h51180636;
temp_data[4043] = 32'h511774a7;
temp_data[4044] = 32'h5116e432;
temp_data[4045] = 32'h511654c5;
temp_data[4046] = 32'h5115c661;
temp_data[4047] = 32'h511538f3;
temp_data[4048] = 32'h5114ac75;
temp_data[4049] = 32'h511420e2;
temp_data[4050] = 32'h5113962d;
temp_data[4051] = 32'h51130c4e;
temp_data[4052] = 32'h51128345;
temp_data[4053] = 32'h5111fb05;
temp_data[4054] = 32'h5111738e;
temp_data[4055] = 32'h5110ecd9;
temp_data[4056] = 32'h511066e0;
temp_data[4057] = 32'h510fe1a0;
temp_data[4058] = 32'h510f5d1c;
temp_data[4059] = 32'h510ed949;
temp_data[4060] = 32'h510e562e;
temp_data[4061] = 32'h510dd3c8;
temp_data[4062] = 32'h510d521a;
temp_data[4063] = 32'h510cd128;
temp_data[4064] = 32'h510c50f4;
temp_data[4065] = 32'h510bd181;
temp_data[4066] = 32'h510b52db;
temp_data[4067] = 32'h510ad50b;
temp_data[4068] = 32'h510a5815;
temp_data[4069] = 32'h5109dc12;
temp_data[4070] = 32'h51096107;
temp_data[4071] = 32'h5108e70c;
temp_data[4072] = 32'h51086e33;
temp_data[4073] = 32'h5107f694;
temp_data[4074] = 32'h51078052;
temp_data[4075] = 32'h51070b85;
temp_data[4076] = 32'h51069852;
temp_data[4077] = 32'h510626e9;
temp_data[4078] = 32'h5105b76f;
temp_data[4079] = 32'h51054a23;
temp_data[4080] = 32'h5104df3b;
temp_data[4081] = 32'h510476fb;
temp_data[4082] = 32'h510411a9;
temp_data[4083] = 32'h5103af9f;
temp_data[4084] = 32'h5103513b;
temp_data[4085] = 32'h5102f6e4;
temp_data[4086] = 32'h5102a112;
temp_data[4087] = 32'h51025048;
temp_data[4088] = 32'h51020518;
temp_data[4089] = 32'h5101c02b;
temp_data[4090] = 32'h51018230;
temp_data[4091] = 32'h51014bfd;
temp_data[4092] = 32'h51011e6d;
temp_data[4093] = 32'h5100fa7f;
temp_data[4094] = 32'h5100e154;
temp_data[4095] = 32'h5100d420;
temp_data[4096] = 32'h50f6dd90;
temp_data[4097] = 32'h50f6e9f7;
temp_data[4098] = 32'h50f7018e;
temp_data[4099] = 32'h50f72325;
temp_data[4100] = 32'h50f74da9;
temp_data[4101] = 32'h50f7801f;
temp_data[4102] = 32'h50f7b9ae;
temp_data[4103] = 32'h50f7f98b;
temp_data[4104] = 32'h50f83f03;
temp_data[4105] = 32'h50f88976;
temp_data[4106] = 32'h50f8d856;
temp_data[4107] = 32'h50f92b1f;
temp_data[4108] = 32'h50f9815e;
temp_data[4109] = 32'h50f9daad;
temp_data[4110] = 32'h50fa36b1;
temp_data[4111] = 32'h50fa9514;
temp_data[4112] = 32'h50faf590;
temp_data[4113] = 32'h50fb57de;
temp_data[4114] = 32'h50fbbbc7;
temp_data[4115] = 32'h50fc2118;
temp_data[4116] = 32'h50fc87a0;
temp_data[4117] = 32'h50fcef35;
temp_data[4118] = 32'h50fd57b4;
temp_data[4119] = 32'h50fdc0f9;
temp_data[4120] = 32'h50fe2aed;
temp_data[4121] = 32'h50fe9574;
temp_data[4122] = 32'h50ff0075;
temp_data[4123] = 32'h50ff6bdf;
temp_data[4124] = 32'h50ffd7a1;
temp_data[4125] = 32'h510043aa;
temp_data[4126] = 32'h5100aff3;
temp_data[4127] = 32'h51011c69;
temp_data[4128] = 32'h51018905;
temp_data[4129] = 32'h5101f5be;
temp_data[4130] = 32'h51026295;
temp_data[4131] = 32'h5102cf78;
temp_data[4132] = 32'h51033c68;
temp_data[4133] = 32'h5103a965;
temp_data[4134] = 32'h51041666;
temp_data[4135] = 32'h5104836f;
temp_data[4136] = 32'h5104f078;
temp_data[4137] = 32'h51055d81;
temp_data[4138] = 32'h5105ca8e;
temp_data[4139] = 32'h5106379b;
temp_data[4140] = 32'h5106a4ad;
temp_data[4141] = 32'h510711be;
temp_data[4142] = 32'h51077ed8;
temp_data[4143] = 32'h5107ebf6;
temp_data[4144] = 32'h5108591d;
temp_data[4145] = 32'h5108c64c;
temp_data[4146] = 32'h51093387;
temp_data[4147] = 32'h5109a0d3;
temp_data[4148] = 32'h510a0e30;
temp_data[4149] = 32'h510a7ba6;
temp_data[4150] = 32'h510ae932;
temp_data[4151] = 32'h510b56d6;
temp_data[4152] = 32'h510bc49c;
temp_data[4153] = 32'h510c3283;
temp_data[4154] = 32'h510ca094;
temp_data[4155] = 32'h510d0ecb;
temp_data[4156] = 32'h510d7d31;
temp_data[4157] = 32'h510debc8;
temp_data[4158] = 32'h510e5a96;
temp_data[4159] = 32'h510ec99f;
temp_data[4160] = 32'h510f38e3;
temp_data[4161] = 32'h510fa86d;
temp_data[4162] = 32'h5110183b;
temp_data[4163] = 32'h51108859;
temp_data[4164] = 32'h5110f8c2;
temp_data[4165] = 32'h51116983;
temp_data[4166] = 32'h5111da9d;
temp_data[4167] = 32'h51124c12;
temp_data[4168] = 32'h5112bdf1;
temp_data[4169] = 32'h51133034;
temp_data[4170] = 32'h5113a2e4;
temp_data[4171] = 32'h51141605;
temp_data[4172] = 32'h511489a4;
temp_data[4173] = 32'h5114fdbd;
temp_data[4174] = 32'h51157258;
temp_data[4175] = 32'h5115e77d;
temp_data[4176] = 32'h51165d31;
temp_data[4177] = 32'h5116d378;
temp_data[4178] = 32'h51174a5a;
temp_data[4179] = 32'h5117c1db;
temp_data[4180] = 32'h51183a08;
temp_data[4181] = 32'h5118b2dd;
temp_data[4182] = 32'h51192c6b;
temp_data[4183] = 32'h5119a6b5;
temp_data[4184] = 32'h511a21c0;
temp_data[4185] = 32'h511a9d95;
temp_data[4186] = 32'h511b1a3b;
temp_data[4187] = 32'h511b97bb;
temp_data[4188] = 32'h511c161e;
temp_data[4189] = 32'h511c956c;
temp_data[4190] = 32'h511d15ad;
temp_data[4191] = 32'h511d96ea;
temp_data[4192] = 32'h511e192f;
temp_data[4193] = 32'h511e9c84;
temp_data[4194] = 32'h511f20f3;
temp_data[4195] = 32'h511fa687;
temp_data[4196] = 32'h51202d49;
temp_data[4197] = 32'h5120b54a;
temp_data[4198] = 32'h51213e92;
temp_data[4199] = 32'h5121c932;
temp_data[4200] = 32'h51225532;
temp_data[4201] = 32'h5122e2a8;
temp_data[4202] = 32'h5123719b;
temp_data[4203] = 32'h51240221;
temp_data[4204] = 32'h51249446;
temp_data[4205] = 32'h5125281c;
temp_data[4206] = 32'h5125bdba;
temp_data[4207] = 32'h51265532;
temp_data[4208] = 32'h5126ee95;
temp_data[4209] = 32'h512789f8;
temp_data[4210] = 32'h51282778;
temp_data[4211] = 32'h5128c72a;
temp_data[4212] = 32'h5129692b;
temp_data[4213] = 32'h512a0d8d;
temp_data[4214] = 32'h512ab474;
temp_data[4215] = 32'h512b5dff;
temp_data[4216] = 32'h512c0a4a;
temp_data[4217] = 32'h512cb97c;
temp_data[4218] = 32'h512d6bb1;
temp_data[4219] = 32'h512e2110;
temp_data[4220] = 32'h512ed9c7;
temp_data[4221] = 32'h512f95fb;
temp_data[4222] = 32'h513055d6;
temp_data[4223] = 32'h51311983;
temp_data[4224] = 32'h5131e137;
temp_data[4225] = 32'h5132ad21;
temp_data[4226] = 32'h51337d74;
temp_data[4227] = 32'h51345265;
temp_data[4228] = 32'h51352c28;
temp_data[4229] = 32'h51360af2;
temp_data[4230] = 32'h5136eefe;
temp_data[4231] = 32'h5137d884;
temp_data[4232] = 32'h5138c7b4;
temp_data[4233] = 32'h5139bccf;
temp_data[4234] = 32'h513ab802;
temp_data[4235] = 32'h513bb97c;
temp_data[4236] = 32'h513cc166;
temp_data[4237] = 32'h513dcfea;
temp_data[4238] = 32'h513ee51d;
temp_data[4239] = 32'h51400115;
temp_data[4240] = 32'h514123d1;
temp_data[4241] = 32'h51424d44;
temp_data[4242] = 32'h51437d46;
temp_data[4243] = 32'h5144b3a2;
temp_data[4244] = 32'h5145f002;
temp_data[4245] = 32'h514731f0;
temp_data[4246] = 32'h514878d5;
temp_data[4247] = 32'h5149c3f8;
temp_data[4248] = 32'h514b1277;
temp_data[4249] = 32'h514c6345;
temp_data[4250] = 32'h514db539;
temp_data[4251] = 32'h514f0703;
temp_data[4252] = 32'h51505736;
temp_data[4253] = 32'h5151a5f4;
temp_data[4254] = 32'h5152f82b;
temp_data[4255] = 32'h51544c5e;
temp_data[4256] = 32'h5155a130;
temp_data[4257] = 32'h5156f566;
temp_data[4258] = 32'h515847e9;
temp_data[4259] = 32'h515997c0;
temp_data[4260] = 32'h515ae426;
temp_data[4261] = 32'h515c2c77;
temp_data[4262] = 32'h515d7033;
temp_data[4263] = 32'h515eaf04;
temp_data[4264] = 32'h515fe8ab;
temp_data[4265] = 32'h51611d0d;
temp_data[4266] = 32'h51624c1f;
temp_data[4267] = 32'h516375ef;
temp_data[4268] = 32'h51649a99;
temp_data[4269] = 32'h5165ba52;
temp_data[4270] = 32'h5166d556;
temp_data[4271] = 32'h5167ebe6;
temp_data[4272] = 32'h5168fe58;
temp_data[4273] = 32'h516a0d02;
temp_data[4274] = 32'h516b1844;
temp_data[4275] = 32'h516c2086;
temp_data[4276] = 32'h516d262d;
temp_data[4277] = 32'h516e29b3;
temp_data[4278] = 32'h516f2b88;
temp_data[4279] = 32'h51702c30;
temp_data[4280] = 32'h51712c28;
temp_data[4281] = 32'h51722bfe;
temp_data[4282] = 32'h51732c3d;
temp_data[4283] = 32'h51742d84;
temp_data[4284] = 32'h51753073;
temp_data[4285] = 32'h517635b5;
temp_data[4286] = 32'h51773e03;
temp_data[4287] = 32'h51784a1f;
temp_data[4288] = 32'h51795ad9;
temp_data[4289] = 32'h517a711d;
temp_data[4290] = 32'h517b8dd6;
temp_data[4291] = 32'h517cb214;
temp_data[4292] = 32'h517ddef8;
temp_data[4293] = 32'h517f15be;
temp_data[4294] = 32'h518057b8;
temp_data[4295] = 32'h5181a66e;
temp_data[4296] = 32'h51830371;
temp_data[4297] = 32'h5184708f;
temp_data[4298] = 32'h5185efbf;
temp_data[4299] = 32'h5187832c;
temp_data[4300] = 32'h51892d34;
temp_data[4301] = 32'h518af080;
temp_data[4302] = 32'h518ccffa;
temp_data[4303] = 32'h518ecee6;
temp_data[4304] = 32'h5190f0d0;
temp_data[4305] = 32'h519339b9;
temp_data[4306] = 32'h5195ae0c;
temp_data[4307] = 32'h519852b5;
temp_data[4308] = 32'h519b2d23;
temp_data[4309] = 32'h519e4367;
temp_data[4310] = 32'h51a19c45;
temp_data[4311] = 32'h51a53f3e;
temp_data[4312] = 32'h51a934a0;
temp_data[4313] = 32'h51ad85be;
temp_data[4314] = 32'h51b23cea;
temp_data[4315] = 32'h51b7659d;
temp_data[4316] = 32'h51bd0ca2;
temp_data[4317] = 32'h51c3401c;
temp_data[4318] = 32'h51ca0fd4;
temp_data[4319] = 32'h51d18d37;
temp_data[4320] = 32'h51d9cb96;
temp_data[4321] = 32'h51e2e054;
temp_data[4322] = 32'h51ece30d;
temp_data[4323] = 32'h51f7edd9;
temp_data[4324] = 32'h52024684;
temp_data[4325] = 32'h520b9247;
temp_data[4326] = 32'h5213e942;
temp_data[4327] = 32'h521b6102;
temp_data[4328] = 32'h52220cb3;
temp_data[4329] = 32'h5227fd44;
temp_data[4330] = 32'h522d419e;
temp_data[4331] = 32'h5231e6bc;
temp_data[4332] = 32'h5235f7cf;
temp_data[4333] = 32'h52397e67;
temp_data[4334] = 32'h523c8273;
temp_data[4335] = 32'h523f0a74;
temp_data[4336] = 32'h52411b7e;
temp_data[4337] = 32'h5242b956;
temp_data[4338] = 32'h5243e671;
temp_data[4339] = 32'h5244a409;
temp_data[4340] = 32'h5244f21b;
temp_data[4341] = 32'h5244cf70;
temp_data[4342] = 32'h5244398f;
temp_data[4343] = 32'h52432cd4;
temp_data[4344] = 32'h5241a448;
temp_data[4345] = 32'h523f99af;
temp_data[4346] = 32'h523d0568;
temp_data[4347] = 32'h5239de72;
temp_data[4348] = 32'h52361a37;
temp_data[4349] = 32'h5231ac93;
temp_data[4350] = 32'h522c8798;
temp_data[4351] = 32'h52269b89;
temp_data[4352] = 32'h521fd677;
temp_data[4353] = 32'h5219f9ec;
temp_data[4354] = 32'h5214f417;
temp_data[4355] = 32'h5210b563;
temp_data[4356] = 32'h520d302f;
temp_data[4357] = 32'h520a58b4;
temp_data[4358] = 32'h520824dd;
temp_data[4359] = 32'h52068c37;
temp_data[4360] = 32'h520587d7;
temp_data[4361] = 32'h5205124d;
temp_data[4362] = 32'h52052795;
temp_data[4363] = 32'h5205c50d;
temp_data[4364] = 32'h5206e979;
temp_data[4365] = 32'h520894f2;
temp_data[4366] = 32'h520ac900;
temp_data[4367] = 32'h520d887f;
temp_data[4368] = 32'h5210d7c3;
temp_data[4369] = 32'h5214bca5;
temp_data[4370] = 32'h52193e81;
temp_data[4371] = 32'h521e6666;
temp_data[4372] = 32'h52243f18;
temp_data[4373] = 32'h522ad545;
temp_data[4374] = 32'h523237a0;
temp_data[4375] = 32'h523a770c;
temp_data[4376] = 32'h5243a6d2;
temp_data[4377] = 32'h524ddcdf;
temp_data[4378] = 32'h525931f9;
temp_data[4379] = 32'h5265c209;
temp_data[4380] = 32'h5273ac7e;
temp_data[4381] = 32'h52831494;
temp_data[4382] = 32'h529421c9;
temp_data[4383] = 32'h52a70047;
temp_data[4384] = 32'h52bbe169;
temp_data[4385] = 32'h52d2fc44;
temp_data[4386] = 32'h52ec8e43;
temp_data[4387] = 32'h5308dbc2;
temp_data[4388] = 32'h532830d7;
temp_data[4389] = 32'h534ae209;
temp_data[4390] = 32'h53714d16;
temp_data[4391] = 32'h539bd9ec;
temp_data[4392] = 32'h53cafb9c;
temp_data[4393] = 32'h53ff3183;
temp_data[4394] = 32'h543474b8;
temp_data[4395] = 32'h54647718;
temp_data[4396] = 32'h548fbab2;
temp_data[4397] = 32'h54b6b4dd;
temp_data[4398] = 32'h54d9cf8d;
temp_data[4399] = 32'h54f96a6a;
temp_data[4400] = 32'h5515dba5;
temp_data[4401] = 32'h552f70c5;
temp_data[4402] = 32'h55466f82;
temp_data[4403] = 32'h555b1666;
temp_data[4404] = 32'h556d9d8c;
temp_data[4405] = 32'h557e3726;
temp_data[4406] = 32'h558d1017;
temp_data[4407] = 32'h559a507a;
temp_data[4408] = 32'h55a61c04;
temp_data[4409] = 32'h55b09281;
temp_data[4410] = 32'h55b9d024;
temp_data[4411] = 32'h55c1edd5;
temp_data[4412] = 32'h55c90193;
temp_data[4413] = 32'h55cf1e9b;
temp_data[4414] = 32'h55d455b4;
temp_data[4415] = 32'h55d8b557;
temp_data[4416] = 32'h55dc49d8;
temp_data[4417] = 32'h55df1d97;
temp_data[4418] = 32'h55e1390d;
temp_data[4419] = 32'h55e2a2f9;
temp_data[4420] = 32'h55e36067;
temp_data[4421] = 32'h55e374c5;
temp_data[4422] = 32'h55e2e1e3;
temp_data[4423] = 32'h55e1a80d;
temp_data[4424] = 32'h55dfc5f4;
temp_data[4425] = 32'h55dd38c1;
temp_data[4426] = 32'h55d9fbf8;
temp_data[4427] = 32'h55d60981;
temp_data[4428] = 32'h55d15986;
temp_data[4429] = 32'h55cbe261;
temp_data[4430] = 32'h55c59885;
temp_data[4431] = 32'h55be6e50;
temp_data[4432] = 32'h55b653f8;
temp_data[4433] = 32'h55ad373f;
temp_data[4434] = 32'h55a30360;
temp_data[4435] = 32'h5597a0b6;
temp_data[4436] = 32'h558af480;
temp_data[4437] = 32'h557ce098;
temp_data[4438] = 32'h556d4313;
temp_data[4439] = 32'h555bf5e0;
temp_data[4440] = 32'h5548ce57;
temp_data[4441] = 32'h55339cbf;
temp_data[4442] = 32'h551c2bd0;
temp_data[4443] = 32'h55023fff;
temp_data[4444] = 32'h54e596ff;
temp_data[4445] = 32'h54c5e6f7;
temp_data[4446] = 32'h54a2ddc2;
temp_data[4447] = 32'h547c2021;
temp_data[4448] = 32'h545148e4;
temp_data[4449] = 32'h5421e7da;
temp_data[4450] = 32'h53ed80e9;
temp_data[4451] = 32'h53b38a65;
temp_data[4452] = 32'h537cecf6;
temp_data[4453] = 32'h534b7968;
temp_data[4454] = 32'h531eae3a;
temp_data[4455] = 32'h52f61659;
temp_data[4456] = 32'h52d14802;
temp_data[4457] = 32'h52afe3ac;
temp_data[4458] = 32'h52919321;
temp_data[4459] = 32'h527608b3;
temp_data[4460] = 32'h525cfe76;
temp_data[4461] = 32'h52463565;
temp_data[4462] = 32'h523174de;
temp_data[4463] = 32'h521e89ec;
temp_data[4464] = 32'h520d46b2;
temp_data[4465] = 32'h51fd8206;
temp_data[4466] = 32'h51ef16ce;
temp_data[4467] = 32'h51e1e3b9;
temp_data[4468] = 32'h51d5cac9;
temp_data[4469] = 32'h51cab10c;
temp_data[4470] = 32'h51c07e35;
temp_data[4471] = 32'h51b71c6d;
temp_data[4472] = 32'h51ae7807;
temp_data[4473] = 32'h51a67f52;
temp_data[4474] = 32'h519f224b;
temp_data[4475] = 32'h51985297;
temp_data[4476] = 32'h5192033a;
temp_data[4477] = 32'h518c2885;
temp_data[4478] = 32'h5186b7e5;
temp_data[4479] = 32'h5181a7d2;
temp_data[4480] = 32'h517cefae;
temp_data[4481] = 32'h517887be;
temp_data[4482] = 32'h517468f1;
temp_data[4483] = 32'h51708cef;
temp_data[4484] = 32'h516cedfe;
temp_data[4485] = 32'h516986e4;
temp_data[4486] = 32'h516652eb;
temp_data[4487] = 32'h51634dd3;
temp_data[4488] = 32'h516073b8;
temp_data[4489] = 32'h515dc11e;
temp_data[4490] = 32'h515b32cf;
temp_data[4491] = 32'h5158c5ef;
temp_data[4492] = 32'h515677d5;
temp_data[4493] = 32'h51544624;
temp_data[4494] = 32'h51522eae;
temp_data[4495] = 32'h51502f77;
temp_data[4496] = 32'h514e46ae;
temp_data[4497] = 32'h514c72b4;
temp_data[4498] = 32'h514ab203;
temp_data[4499] = 32'h51490343;
temp_data[4500] = 32'h51476530;
temp_data[4501] = 32'h5145d6a1;
temp_data[4502] = 32'h51445693;
temp_data[4503] = 32'h5142e404;
temp_data[4504] = 32'h51417e17;
temp_data[4505] = 32'h514023ff;
temp_data[4506] = 32'h513ed4f6;
temp_data[4507] = 32'h513d9058;
temp_data[4508] = 32'h513c5575;
temp_data[4509] = 32'h513b23c4;
temp_data[4510] = 32'h5139fab5;
temp_data[4511] = 32'h5138d9cb;
temp_data[4512] = 32'h5137c090;
temp_data[4513] = 32'h5136ae97;
temp_data[4514] = 32'h5135a377;
temp_data[4515] = 32'h51349ed8;
temp_data[4516] = 32'h5133a05e;
temp_data[4517] = 32'h5132a7b5;
temp_data[4518] = 32'h5131b49a;
temp_data[4519] = 32'h5130c6bd;
temp_data[4520] = 32'h512fdde3;
temp_data[4521] = 32'h512ef9ca;
temp_data[4522] = 32'h512e1a37;
temp_data[4523] = 32'h512d3ef7;
temp_data[4524] = 32'h512c67d7;
temp_data[4525] = 32'h512b94a3;
temp_data[4526] = 32'h512ac52e;
temp_data[4527] = 32'h5129f951;
temp_data[4528] = 32'h512930e4;
temp_data[4529] = 32'h51286bba;
temp_data[4530] = 32'h5127a9b5;
temp_data[4531] = 32'h5126eab3;
temp_data[4532] = 32'h51262e90;
temp_data[4533] = 32'h51257532;
temp_data[4534] = 32'h5124be77;
temp_data[4535] = 32'h51240a46;
temp_data[4536] = 32'h51235882;
temp_data[4537] = 32'h5122a915;
temp_data[4538] = 32'h5121fbe7;
temp_data[4539] = 32'h512150df;
temp_data[4540] = 32'h5120a7e7;
temp_data[4541] = 32'h512000eb;
temp_data[4542] = 32'h511f5bd5;
temp_data[4543] = 32'h511eb899;
temp_data[4544] = 32'h511e171a;
temp_data[4545] = 32'h511d774b;
temp_data[4546] = 32'h511cd91f;
temp_data[4547] = 32'h511c3c82;
temp_data[4548] = 32'h511ba162;
temp_data[4549] = 32'h511b07b8;
temp_data[4550] = 32'h511a6f69;
temp_data[4551] = 32'h5119d873;
temp_data[4552] = 32'h511942c8;
temp_data[4553] = 32'h5118ae53;
temp_data[4554] = 32'h51181b0d;
temp_data[4555] = 32'h511788ec;
temp_data[4556] = 32'h5116f7e4;
temp_data[4557] = 32'h511667e8;
temp_data[4558] = 32'h5115d8f1;
temp_data[4559] = 32'h51154af5;
temp_data[4560] = 32'h5114bde8;
temp_data[4561] = 32'h511431c6;
temp_data[4562] = 32'h5113a683;
temp_data[4563] = 32'h51131c1d;
temp_data[4564] = 32'h51129286;
temp_data[4565] = 32'h511209c0;
temp_data[4566] = 32'h511181bf;
temp_data[4567] = 32'h5110fa7f;
temp_data[4568] = 32'h51107400;
temp_data[4569] = 32'h510fee3d;
temp_data[4570] = 32'h510f6934;
temp_data[4571] = 32'h510ee4de;
temp_data[4572] = 32'h510e6141;
temp_data[4573] = 32'h510dde59;
temp_data[4574] = 32'h510d5c2d;
temp_data[4575] = 32'h510cdaba;
temp_data[4576] = 32'h510c5a08;
temp_data[4577] = 32'h510bda1b;
temp_data[4578] = 32'h510b5afb;
temp_data[4579] = 32'h510adcad;
temp_data[4580] = 32'h510a5f46;
temp_data[4581] = 32'h5109e2ca;
temp_data[4582] = 32'h51096749;
temp_data[4583] = 32'h5108ecd9;
temp_data[4584] = 32'h51087393;
temp_data[4585] = 32'h5107fb87;
temp_data[4586] = 32'h510784d3;
temp_data[4587] = 32'h51070f9d;
temp_data[4588] = 32'h51069c02;
temp_data[4589] = 32'h51062a35;
temp_data[4590] = 32'h5105ba5a;
temp_data[4591] = 32'h51054cad;
temp_data[4592] = 32'h5104e165;
temp_data[4593] = 32'h510478cd;
temp_data[4594] = 32'h51041327;
temp_data[4595] = 32'h5103b0c9;
temp_data[4596] = 32'h5103521a;
temp_data[4597] = 32'h5102f777;
temp_data[4598] = 32'h5102a162;
temp_data[4599] = 32'h51025059;
temp_data[4600] = 32'h510204ee;
temp_data[4601] = 32'h5101bfcf;
temp_data[4602] = 32'h510181a6;
temp_data[4603] = 32'h51014b49;
temp_data[4604] = 32'h51011d9b;
temp_data[4605] = 32'h5100f99c;
temp_data[4606] = 32'h5100e05d;
temp_data[4607] = 32'h5100d320;
temp_data[4608] = 32'h50f6d1bf;
temp_data[4609] = 32'h50f6de2b;
temp_data[4610] = 32'h50f6f5cf;
temp_data[4611] = 32'h50f71776;
temp_data[4612] = 32'h50f7420f;
temp_data[4613] = 32'h50f774a3;
temp_data[4614] = 32'h50f7ae58;
temp_data[4615] = 32'h50f7ee5b;
temp_data[4616] = 32'h50f83401;
temp_data[4617] = 32'h50f87eaa;
temp_data[4618] = 32'h50f8cdc0;
temp_data[4619] = 32'h50f920c9;
temp_data[4620] = 32'h50f9774b;
temp_data[4621] = 32'h50f9d0dd;
temp_data[4622] = 32'h50fa2d2c;
temp_data[4623] = 32'h50fa8bdf;
temp_data[4624] = 32'h50faeca7;
temp_data[4625] = 32'h50fb4f4c;
temp_data[4626] = 32'h50fbb38d;
temp_data[4627] = 32'h50fc1937;
temp_data[4628] = 32'h50fc8017;
temp_data[4629] = 32'h50fce80c;
temp_data[4630] = 32'h50fd50ec;
temp_data[4631] = 32'h50fdba95;
temp_data[4632] = 32'h50fe24ee;
temp_data[4633] = 32'h50fe8fda;
temp_data[4634] = 32'h50fefb44;
temp_data[4635] = 32'h50ff671b;
temp_data[4636] = 32'h50ffd346;
temp_data[4637] = 32'h51003fc0;
temp_data[4638] = 32'h5100ac71;
temp_data[4639] = 32'h51011959;
temp_data[4640] = 32'h51018666;
temp_data[4641] = 32'h5101f395;
temp_data[4642] = 32'h510260d9;
temp_data[4643] = 32'h5102ce31;
temp_data[4644] = 32'h51033b9b;
temp_data[4645] = 32'h5103a90d;
temp_data[4646] = 32'h51041683;
temp_data[4647] = 32'h51048402;
temp_data[4648] = 32'h5104f184;
temp_data[4649] = 32'h51055f07;
temp_data[4650] = 32'h5105cc8e;
temp_data[4651] = 32'h51063a19;
temp_data[4652] = 32'h5106a7a4;
temp_data[4653] = 32'h51071533;
temp_data[4654] = 32'h510782cb;
temp_data[4655] = 32'h5107f067;
temp_data[4656] = 32'h51085e0b;
temp_data[4657] = 32'h5108cbbc;
temp_data[4658] = 32'h5109397a;
temp_data[4659] = 32'h5109a748;
temp_data[4660] = 32'h510a1527;
temp_data[4661] = 32'h510a831b;
temp_data[4662] = 32'h510af12c;
temp_data[4663] = 32'h510b5f57;
temp_data[4664] = 32'h510bcda3;
temp_data[4665] = 32'h510c3c10;
temp_data[4666] = 32'h510caaa4;
temp_data[4667] = 32'h510d1965;
temp_data[4668] = 32'h510d8851;
temp_data[4669] = 32'h510df773;
temp_data[4670] = 32'h510e66cb;
temp_data[4671] = 32'h510ed65e;
temp_data[4672] = 32'h510f4630;
temp_data[4673] = 32'h510fb646;
temp_data[4674] = 32'h511026a2;
temp_data[4675] = 32'h5110974a;
temp_data[4676] = 32'h51110846;
temp_data[4677] = 32'h51117996;
temp_data[4678] = 32'h5111eb42;
temp_data[4679] = 32'h51125d4a;
temp_data[4680] = 32'h5112cfbc;
temp_data[4681] = 32'h51134291;
temp_data[4682] = 32'h5113b5d9;
temp_data[4683] = 32'h51142995;
temp_data[4684] = 32'h51149dc7;
temp_data[4685] = 32'h5115127b;
temp_data[4686] = 32'h511587b1;
temp_data[4687] = 32'h5115fd72;
temp_data[4688] = 32'h511673c5;
temp_data[4689] = 32'h5116eaab;
temp_data[4690] = 32'h5117622c;
temp_data[4691] = 32'h5117da55;
temp_data[4692] = 32'h51185322;
temp_data[4693] = 32'h5118cc9f;
temp_data[4694] = 32'h511946d4;
temp_data[4695] = 32'h5119c1c6;
temp_data[4696] = 32'h511a3d7d;
temp_data[4697] = 32'h511aba02;
temp_data[4698] = 32'h511b3758;
temp_data[4699] = 32'h511bb58d;
temp_data[4700] = 32'h511c34a4;
temp_data[4701] = 32'h511cb4ab;
temp_data[4702] = 32'h511d35a4;
temp_data[4703] = 32'h511db7a2;
temp_data[4704] = 32'h511e3aa3;
temp_data[4705] = 32'h511ebeba;
temp_data[4706] = 32'h511f43f2;
temp_data[4707] = 32'h511fca4f;
temp_data[4708] = 32'h512051e3;
temp_data[4709] = 32'h5120dab6;
temp_data[4710] = 32'h512164d4;
temp_data[4711] = 32'h5121f052;
temp_data[4712] = 32'h51227d35;
temp_data[4713] = 32'h51230b8d;
temp_data[4714] = 32'h51239b6f;
temp_data[4715] = 32'h51242ce9;
temp_data[4716] = 32'h5124c005;
temp_data[4717] = 32'h512554de;
temp_data[4718] = 32'h5125eb89;
temp_data[4719] = 32'h51268412;
temp_data[4720] = 32'h51271e93;
temp_data[4721] = 32'h5127bb1f;
temp_data[4722] = 32'h512859d1;
temp_data[4723] = 32'h5128fac2;
temp_data[4724] = 32'h51299e0e;
temp_data[4725] = 32'h512a43d0;
temp_data[4726] = 32'h512aec25;
temp_data[4727] = 32'h512b9731;
temp_data[4728] = 32'h512c450f;
temp_data[4729] = 32'h512cf5ed;
temp_data[4730] = 32'h512da9e7;
temp_data[4731] = 32'h512e6128;
temp_data[4732] = 32'h512f1bdf;
temp_data[4733] = 32'h512fda30;
temp_data[4734] = 32'h51309c52;
temp_data[4735] = 32'h5131626f;
temp_data[4736] = 32'h51322cc3;
temp_data[4737] = 32'h5132fb7f;
temp_data[4738] = 32'h5133cedd;
temp_data[4739] = 32'h5134a716;
temp_data[4740] = 32'h51358466;
temp_data[4741] = 32'h5136670e;
temp_data[4742] = 32'h51374f4c;
temp_data[4743] = 32'h51383d64;
temp_data[4744] = 32'h51393194;
temp_data[4745] = 32'h513a2c1f;
temp_data[4746] = 32'h513b2d41;
temp_data[4747] = 32'h513c3537;
temp_data[4748] = 32'h513d4439;
temp_data[4749] = 32'h513e5a79;
temp_data[4750] = 32'h513f7825;
temp_data[4751] = 32'h51409d56;
temp_data[4752] = 32'h5141ca21;
temp_data[4753] = 32'h5142fe82;
temp_data[4754] = 32'h51443a64;
temp_data[4755] = 32'h51457d9a;
temp_data[4756] = 32'h5146c7d2;
temp_data[4757] = 32'h5148189c;
temp_data[4758] = 32'h51496f5d;
temp_data[4759] = 32'h514acb4f;
temp_data[4760] = 32'h514c2b80;
temp_data[4761] = 32'h514d8ece;
temp_data[4762] = 32'h514ef3e4;
temp_data[4763] = 32'h5150594b;
temp_data[4764] = 32'h5151bd62;
temp_data[4765] = 32'h51532014;
temp_data[4766] = 32'h51548612;
temp_data[4767] = 32'h5155edb3;
temp_data[4768] = 32'h51575565;
temp_data[4769] = 32'h5158bbc3;
temp_data[4770] = 32'h515a1f92;
temp_data[4771] = 32'h515b7fcc;
temp_data[4772] = 32'h515cdb90;
temp_data[4773] = 32'h515e3240;
temp_data[4774] = 32'h515f8356;
temp_data[4775] = 32'h5160ce7d;
temp_data[4776] = 32'h51621383;
temp_data[4777] = 32'h51635254;
temp_data[4778] = 32'h51648af8;
temp_data[4779] = 32'h5165bd84;
temp_data[4780] = 32'h5166ea2d;
temp_data[4781] = 32'h5168112c;
temp_data[4782] = 32'h516932ca;
temp_data[4783] = 32'h516a4f5d;
temp_data[4784] = 32'h516b6745;
temp_data[4785] = 32'h516c7ae1;
temp_data[4786] = 32'h516d8aa0;
temp_data[4787] = 32'h516e96ee;
temp_data[4788] = 32'h516fa045;
temp_data[4789] = 32'h5170a716;
temp_data[4790] = 32'h5171abe7;
temp_data[4791] = 32'h5172af3a;
temp_data[4792] = 32'h5173b196;
temp_data[4793] = 32'h5174b38d;
temp_data[4794] = 32'h5175b5af;
temp_data[4795] = 32'h5176b895;
temp_data[4796] = 32'h5177bced;
temp_data[4797] = 32'h5178c361;
temp_data[4798] = 32'h5179cca7;
temp_data[4799] = 32'h517ad988;
temp_data[4800] = 32'h517bead5;
temp_data[4801] = 32'h517d0171;
temp_data[4802] = 32'h517e1e54;
temp_data[4803] = 32'h517f4281;
temp_data[4804] = 32'h51806f1a;
temp_data[4805] = 32'h5181a555;
temp_data[4806] = 32'h5182e68e;
temp_data[4807] = 32'h5184343b;
temp_data[4808] = 32'h51858ff3;
temp_data[4809] = 32'h5186fb7a;
temp_data[4810] = 32'h518878c0;
temp_data[4811] = 32'h518a09ea;
temp_data[4812] = 32'h518bb153;
temp_data[4813] = 32'h518d719b;
temp_data[4814] = 32'h518f4da1;
temp_data[4815] = 32'h51914899;
temp_data[4816] = 32'h51936613;
temp_data[4817] = 32'h5195aa00;
temp_data[4818] = 32'h519818b9;
temp_data[4819] = 32'h519ab720;
temp_data[4820] = 32'h519d8a98;
temp_data[4821] = 32'h51a0992d;
temp_data[4822] = 32'h51a3e985;
temp_data[4823] = 32'h51a7831f;
temp_data[4824] = 32'h51ab6e44;
temp_data[4825] = 32'h51afb431;
temp_data[4826] = 32'h51b45f39;
temp_data[4827] = 32'h51b97ad5;
temp_data[4828] = 32'h51bf13cb;
temp_data[4829] = 32'h51c53850;
temp_data[4830] = 32'h51cbf83c;
temp_data[4831] = 32'h51d36517;
temp_data[4832] = 32'h51db9258;
temp_data[4833] = 32'h51e4958e;
temp_data[4834] = 32'h51ee867f;
temp_data[4835] = 32'h51f97f8d;
temp_data[4836] = 32'h5203c6b5;
temp_data[4837] = 32'h520d016d;
temp_data[4838] = 32'h5215480f;
temp_data[4839] = 32'h521cb04f;
temp_data[4840] = 32'h52234d83;
temp_data[4841] = 32'h522930be;
temp_data[4842] = 32'h522e68f9;
temp_data[4843] = 32'h5233033e;
temp_data[4844] = 32'h52370abf;
temp_data[4845] = 32'h523a890d;
temp_data[4846] = 32'h523d860e;
temp_data[4847] = 32'h5240083a;
temp_data[4848] = 32'h5242149c;
temp_data[4849] = 32'h5243aee6;
temp_data[4850] = 32'h5244d97f;
temp_data[4851] = 32'h52459592;
temp_data[4852] = 32'h5245e300;
temp_data[4853] = 32'h5245c087;
temp_data[4854] = 32'h52452ba1;
temp_data[4855] = 32'h5244208e;
temp_data[4856] = 32'h52429a46;
temp_data[4857] = 32'h52409279;
temp_data[4858] = 32'h523e017e;
temp_data[4859] = 32'h523ade2f;
temp_data[4860] = 32'h52371df7;
temp_data[4861] = 32'h5232b491;
temp_data[4862] = 32'h522d9403;
temp_data[4863] = 32'h5227ac75;
temp_data[4864] = 32'h5220ebf6;
temp_data[4865] = 32'h521b13e8;
temp_data[4866] = 32'h52161277;
temp_data[4867] = 32'h5211d7f5;
temp_data[4868] = 32'h520e56ac;
temp_data[4869] = 32'h520b82c3;
temp_data[4870] = 32'h5209520d;
temp_data[4871] = 32'h5207bc0a;
temp_data[4872] = 32'h5206b9b6;
temp_data[4873] = 32'h52064591;
temp_data[4874] = 32'h52065b79;
temp_data[4875] = 32'h5206f8ba;
temp_data[4876] = 32'h52081c00;
temp_data[4877] = 32'h5209c554;
temp_data[4878] = 32'h520bf612;
temp_data[4879] = 32'h520eb103;
temp_data[4880] = 32'h5211fa66;
temp_data[4881] = 32'h5215d7e9;
temp_data[4882] = 32'h521a50ca;
temp_data[4883] = 32'h521f6df0;
temp_data[4884] = 32'h52253a00;
temp_data[4885] = 32'h522bc172;
temp_data[4886] = 32'h523312d3;
temp_data[4887] = 32'h523b3ed5;
temp_data[4888] = 32'h5244588e;
temp_data[4889] = 32'h524e75b0;
temp_data[4890] = 32'h5259aec9;
temp_data[4891] = 32'h52661f8e;
temp_data[4892] = 32'h5273e732;
temp_data[4893] = 32'h528328b7;
temp_data[4894] = 32'h52940b63;
temp_data[4895] = 32'h52a6bb38;
temp_data[4896] = 32'h52bb696e;
temp_data[4897] = 32'h52d24cfd;
temp_data[4898] = 32'h52eba351;
temp_data[4899] = 32'h5307b0e2;
temp_data[4900] = 32'h5326c1f0;
temp_data[4901] = 32'h53492b5a;
temp_data[4902] = 32'h536f4b5e;
temp_data[4903] = 32'h53998a83;
temp_data[4904] = 32'h53c85c92;
temp_data[4905] = 32'h53fc41c8;
temp_data[4906] = 32'h54313426;
temp_data[4907] = 32'h5460e66d;
temp_data[4908] = 32'h548bdb83;
temp_data[4909] = 32'h54b28987;
temp_data[4910] = 32'h54d55b1d;
temp_data[4911] = 32'h54f4b060;
temp_data[4912] = 32'h5510dfdf;
temp_data[4913] = 32'h552a3761;
temp_data[4914] = 32'h5540fcb9;
temp_data[4915] = 32'h55556e72;
temp_data[4916] = 32'h5567c48f;
temp_data[4917] = 32'h5578312b;
temp_data[4918] = 32'h5586e100;
temp_data[4919] = 32'h5593fbec;
temp_data[4920] = 32'h559fa576;
temp_data[4921] = 32'h55a9fd2f;
temp_data[4922] = 32'h55b31f10;
temp_data[4923] = 32'h55bb23d9;
temp_data[4924] = 32'h55c22147;
temp_data[4925] = 32'h55c82a73;
temp_data[4926] = 32'h55cd4ff0;
temp_data[4927] = 32'h55d1a017;
temp_data[4928] = 32'h55d52718;
temp_data[4929] = 32'h55d7ef31;
temp_data[4930] = 32'h55da00c5;
temp_data[4931] = 32'h55db6280;
temp_data[4932] = 32'h55dc195d;
temp_data[4933] = 32'h55dc28b7;
temp_data[4934] = 32'h55db9260;
temp_data[4935] = 32'h55da5697;
temp_data[4936] = 32'h55d87415;
temp_data[4937] = 32'h55d5e804;
temp_data[4938] = 32'h55d2adf3;
temp_data[4939] = 32'h55cebfdb;
temp_data[4940] = 32'h55ca15f9;
temp_data[4941] = 32'h55c4a6bd;
temp_data[4942] = 32'h55be66b2;
temp_data[4943] = 32'h55b7485e;
temp_data[4944] = 32'h55af3c15;
temp_data[4945] = 32'h55a62fcf;
temp_data[4946] = 32'h559c0ee9;
temp_data[4947] = 32'h5590c1f4;
temp_data[4948] = 32'h55842e6a;
temp_data[4949] = 32'h55763659;
temp_data[4950] = 32'h5566b80b;
temp_data[4951] = 32'h55558da4;
temp_data[4952] = 32'h55428cb0;
temp_data[4953] = 32'h552d85a9;
temp_data[4954] = 32'h5516435f;
temp_data[4955] = 32'h54fc8a5d;
temp_data[4956] = 32'h54e01855;
temp_data[4957] = 32'h54c0a348;
temp_data[4958] = 32'h549dd8dc;
temp_data[4959] = 32'h54775d79;
temp_data[4960] = 32'h544ccb5c;
temp_data[4961] = 32'h541db1c0;
temp_data[4962] = 32'h53e993bc;
temp_data[4963] = 32'h53afe6c9;
temp_data[4964] = 32'h537992b8;
temp_data[4965] = 32'h5348676a;
temp_data[4966] = 32'h531be293;
temp_data[4967] = 32'h52f38e7a;
temp_data[4968] = 32'h52cf00bd;
temp_data[4969] = 32'h52add966;
temp_data[4970] = 32'h528fc209;
temp_data[4971] = 32'h52746cc6;
temp_data[4972] = 32'h525b939f;
temp_data[4973] = 32'h5244f7a9;
temp_data[4974] = 32'h52306057;
temp_data[4975] = 32'h521d9add;
temp_data[4976] = 32'h520c799e;
temp_data[4977] = 32'h51fcd399;
temp_data[4978] = 32'h51ee83fd;
temp_data[4979] = 32'h51e169b1;
temp_data[4980] = 32'h51d566f5;
temp_data[4981] = 32'h51ca610b;
temp_data[4982] = 32'h51c03fdd;
temp_data[4983] = 32'h51b6edd0;
temp_data[4984] = 32'h51ae5764;
temp_data[4985] = 32'h51a66b09;
temp_data[4986] = 32'h519f18f4;
temp_data[4987] = 32'h519852eb;
temp_data[4988] = 32'h51920c0f;
temp_data[4989] = 32'h518c38d2;
temp_data[4990] = 32'h5186cec0;
temp_data[4991] = 32'h5181c469;
temp_data[4992] = 32'h517d1149;
temp_data[4993] = 32'h5178adb0;
temp_data[4994] = 32'h517492a7;
temp_data[4995] = 32'h5170b9e5;
temp_data[4996] = 32'h516d1db8;
temp_data[4997] = 32'h5169b8fe;
temp_data[4998] = 32'h51668705;
temp_data[4999] = 32'h51638399;    
    end
    

initial begin
power_data[0] = 32'h00000086;
power_data[1] = 32'h00000086;
power_data[2] = 32'h00000086;
power_data[3] = 32'h00000086;
power_data[4] = 32'h00000086;
power_data[5] = 32'h00000086;
power_data[6] = 32'h00000086;
power_data[7] = 32'h00000086;
power_data[8] = 32'h00000086;
power_data[9] = 32'h00000086;
power_data[10] = 32'h00000086;
power_data[11] = 32'h00000086;
power_data[12] = 32'h00000086;
power_data[13] = 32'h00000086;
power_data[14] = 32'h00000086;
power_data[15] = 32'h00000086;
power_data[16] = 32'h00000086;
power_data[17] = 32'h00000086;
power_data[18] = 32'h00000086;
power_data[19] = 32'h00000086;
power_data[20] = 32'h00000086;
power_data[21] = 32'h00000086;
power_data[22] = 32'h00000086;
power_data[23] = 32'h00000086;
power_data[24] = 32'h00000086;
power_data[25] = 32'h00000086;
power_data[26] = 32'h00000086;
power_data[27] = 32'h00000086;
power_data[28] = 32'h00000086;
power_data[29] = 32'h00000086;
power_data[30] = 32'h00000086;
power_data[31] = 32'h00000086;
power_data[32] = 32'h00000086;
power_data[33] = 32'h00000086;
power_data[34] = 32'h00000086;
power_data[35] = 32'h00000086;
power_data[36] = 32'h00000086;
power_data[37] = 32'h00000086;
power_data[38] = 32'h00000086;
power_data[39] = 32'h00000086;
power_data[40] = 32'h00000086;
power_data[41] = 32'h00000086;
power_data[42] = 32'h00000086;
power_data[43] = 32'h00000086;
power_data[44] = 32'h00000086;
power_data[45] = 32'h00000086;
power_data[46] = 32'h00000086;
power_data[47] = 32'h00000086;
power_data[48] = 32'h00000086;
power_data[49] = 32'h00000086;
power_data[50] = 32'h00000086;
power_data[51] = 32'h00000086;
power_data[52] = 32'h00000086;
power_data[53] = 32'h00000086;
power_data[54] = 32'h00000086;
power_data[55] = 32'h00000086;
power_data[56] = 32'h00000086;
power_data[57] = 32'h00000086;
power_data[58] = 32'h00000086;
power_data[59] = 32'h00000086;
power_data[60] = 32'h00000086;
power_data[61] = 32'h00000086;
power_data[62] = 32'h00000086;
power_data[63] = 32'h00000086;
power_data[64] = 32'h00000086;
power_data[65] = 32'h00000086;
power_data[66] = 32'h00000086;
power_data[67] = 32'h00000086;
power_data[68] = 32'h00000086;
power_data[69] = 32'h00000086;
power_data[70] = 32'h00000086;
power_data[71] = 32'h00000086;
power_data[72] = 32'h00000086;
power_data[73] = 32'h00000086;
power_data[74] = 32'h00000086;
power_data[75] = 32'h00000086;
power_data[76] = 32'h00000086;
power_data[77] = 32'h00000086;
power_data[78] = 32'h00000086;
power_data[79] = 32'h00000086;
power_data[80] = 32'h00000086;
power_data[81] = 32'h00000086;
power_data[82] = 32'h00000086;
power_data[83] = 32'h00000086;
power_data[84] = 32'h00000086;
power_data[85] = 32'h00000086;
power_data[86] = 32'h00000086;
power_data[87] = 32'h00000086;
power_data[88] = 32'h00000086;
power_data[89] = 32'h00000086;
power_data[90] = 32'h00000086;
power_data[91] = 32'h00000086;
power_data[92] = 32'h00000086;
power_data[93] = 32'h00000086;
power_data[94] = 32'h00000086;
power_data[95] = 32'h00000086;
power_data[96] = 32'h00000086;
power_data[97] = 32'h00000086;
power_data[98] = 32'h00000086;
power_data[99] = 32'h00000086;
power_data[100] = 32'h00000086;
power_data[101] = 32'h00000086;
power_data[102] = 32'h00000086;
power_data[103] = 32'h00000086;
power_data[104] = 32'h00000086;
power_data[105] = 32'h00000086;
power_data[106] = 32'h00000086;
power_data[107] = 32'h00000086;
power_data[108] = 32'h00000086;
power_data[109] = 32'h00000086;
power_data[110] = 32'h00000086;
power_data[111] = 32'h00000086;
power_data[112] = 32'h00000086;
power_data[113] = 32'h00000086;
power_data[114] = 32'h00000086;
power_data[115] = 32'h00000086;
power_data[116] = 32'h00000086;
power_data[117] = 32'h00000086;
power_data[118] = 32'h00000086;
power_data[119] = 32'h00000086;
power_data[120] = 32'h00000086;
power_data[121] = 32'h00000086;
power_data[122] = 32'h00000086;
power_data[123] = 32'h00000086;
power_data[124] = 32'h00000086;
power_data[125] = 32'h00000086;
power_data[126] = 32'h00000086;
power_data[127] = 32'h00000086;
power_data[128] = 32'h00000086;
power_data[129] = 32'h00000086;
power_data[130] = 32'h00000086;
power_data[131] = 32'h00000086;
power_data[132] = 32'h00000086;
power_data[133] = 32'h00000086;
power_data[134] = 32'h00000086;
power_data[135] = 32'h00000086;
power_data[136] = 32'h00000086;
power_data[137] = 32'h00000086;
power_data[138] = 32'h00000086;
power_data[139] = 32'h00000086;
power_data[140] = 32'h00000086;
power_data[141] = 32'h00000086;
power_data[142] = 32'h00000086;
power_data[143] = 32'h00000086;
power_data[144] = 32'h00000086;
power_data[145] = 32'h00000086;
power_data[146] = 32'h00000086;
power_data[147] = 32'h00000086;
power_data[148] = 32'h00000086;
power_data[149] = 32'h00000086;
power_data[150] = 32'h00000086;
power_data[151] = 32'h00000086;
power_data[152] = 32'h00000086;
power_data[153] = 32'h00000086;
power_data[154] = 32'h00000086;
power_data[155] = 32'h00000082;
power_data[156] = 32'h00000069;
power_data[157] = 32'h00000069;
power_data[158] = 32'h00000069;
power_data[159] = 32'h00000069;
power_data[160] = 32'h00000069;
power_data[161] = 32'h00000069;
power_data[162] = 32'h00000069;
power_data[163] = 32'h00000069;
power_data[164] = 32'h00000069;
power_data[165] = 32'h00000069;
power_data[166] = 32'h00000069;
power_data[167] = 32'h00000069;
power_data[168] = 32'h00000069;
power_data[169] = 32'h00000069;
power_data[170] = 32'h00000069;
power_data[171] = 32'h00000069;
power_data[172] = 32'h00000069;
power_data[173] = 32'h00000069;
power_data[174] = 32'h00000069;
power_data[175] = 32'h00000069;
power_data[176] = 32'h00000069;
power_data[177] = 32'h00000069;
power_data[178] = 32'h00000069;
power_data[179] = 32'h00000069;
power_data[180] = 32'h00000069;
power_data[181] = 32'h00000069;
power_data[182] = 32'h00000069;
power_data[183] = 32'h00000069;
power_data[184] = 32'h00000069;
power_data[185] = 32'h00000069;
power_data[186] = 32'h00000069;
power_data[187] = 32'h00000069;
power_data[188] = 32'h00000069;
power_data[189] = 32'h00000069;
power_data[190] = 32'h00000069;
power_data[191] = 32'h00000069;
power_data[192] = 32'h00000069;
power_data[193] = 32'h00000069;
power_data[194] = 32'h00000069;
power_data[195] = 32'h00000069;
power_data[196] = 32'h00000069;
power_data[197] = 32'h00000069;
power_data[198] = 32'h00000069;
power_data[199] = 32'h00000069;
power_data[200] = 32'h00000069;
power_data[201] = 32'h00000069;
power_data[202] = 32'h00000069;
power_data[203] = 32'h00000069;
power_data[204] = 32'h00000069;
power_data[205] = 32'h00000069;
power_data[206] = 32'h00000069;
power_data[207] = 32'h00000069;
power_data[208] = 32'h00000069;
power_data[209] = 32'h00000069;
power_data[210] = 32'h00000069;
power_data[211] = 32'h00000069;
power_data[212] = 32'h00000069;
power_data[213] = 32'h00000069;
power_data[214] = 32'h00000069;
power_data[215] = 32'h00000069;
power_data[216] = 32'h00000069;
power_data[217] = 32'h00000069;
power_data[218] = 32'h00000069;
power_data[219] = 32'h00000069;
power_data[220] = 32'h00000069;
power_data[221] = 32'h00000069;
power_data[222] = 32'h00000069;
power_data[223] = 32'h00000069;
power_data[224] = 32'h00000069;
power_data[225] = 32'h00000069;
power_data[226] = 32'h0000077d;
power_data[227] = 32'h00000942;
power_data[228] = 32'h00000942;
power_data[229] = 32'h00000942;
power_data[230] = 32'h00000942;
power_data[231] = 32'h00000942;
power_data[232] = 32'h00000942;
power_data[233] = 32'h00000942;
power_data[234] = 32'h00000942;
power_data[235] = 32'h00000942;
power_data[236] = 32'h00000942;
power_data[237] = 32'h00000942;
power_data[238] = 32'h00000942;
power_data[239] = 32'h00000942;
power_data[240] = 32'h00000942;
power_data[241] = 32'h00000942;
power_data[242] = 32'h00000942;
power_data[243] = 32'h00000942;
power_data[244] = 32'h00000942;
power_data[245] = 32'h00000942;
power_data[246] = 32'h00000942;
power_data[247] = 32'h00000942;
power_data[248] = 32'h00000942;
power_data[249] = 32'h00000942;
power_data[250] = 32'h00000942;
power_data[251] = 32'h00000942;
power_data[252] = 32'h00000942;
power_data[253] = 32'h00000942;
power_data[254] = 32'h00000942;
power_data[255] = 32'h00000232;
power_data[256] = 32'h00000232;
power_data[257] = 32'h00000232;
power_data[258] = 32'h00000232;
power_data[259] = 32'h00000232;
power_data[260] = 32'h00000232;
power_data[261] = 32'h00000232;
power_data[262] = 32'h00000232;
power_data[263] = 32'h00000232;
power_data[264] = 32'h00000232;
power_data[265] = 32'h00000232;
power_data[266] = 32'h00000232;
power_data[267] = 32'h00000232;
power_data[268] = 32'h00000232;
power_data[269] = 32'h00000232;
power_data[270] = 32'h00000232;
power_data[271] = 32'h00000232;
power_data[272] = 32'h00000232;
power_data[273] = 32'h00000232;
power_data[274] = 32'h00000232;
power_data[275] = 32'h00000232;
power_data[276] = 32'h00000232;
power_data[277] = 32'h00000232;
power_data[278] = 32'h00000232;
power_data[279] = 32'h00000232;
power_data[280] = 32'h00000232;
power_data[281] = 32'h00000232;
power_data[282] = 32'h00000232;
power_data[283] = 32'h00000232;
power_data[284] = 32'h00000232;
power_data[285] = 32'h00000232;
power_data[286] = 32'h00000232;
power_data[287] = 32'h00000232;
power_data[288] = 32'h00000232;
power_data[289] = 32'h00000232;
power_data[290] = 32'h00000232;
power_data[291] = 32'h00000232;
power_data[292] = 32'h00000232;
power_data[293] = 32'h00000232;
power_data[294] = 32'h00000232;
power_data[295] = 32'h00000232;
power_data[296] = 32'h000013d3;
power_data[297] = 32'h00002e41;
power_data[298] = 32'h00002e41;
power_data[299] = 32'h00002e41;
power_data[300] = 32'h00002e41;
power_data[301] = 32'h00002e41;
power_data[302] = 32'h00002e41;
power_data[303] = 32'h00002e41;
power_data[304] = 32'h00002e41;
power_data[305] = 32'h00002e41;
power_data[306] = 32'h00002e41;
power_data[307] = 32'h00002e41;
power_data[308] = 32'h00002e41;
power_data[309] = 32'h00002e41;
power_data[310] = 32'h00002e41;
power_data[311] = 32'h00002e41;
power_data[312] = 32'h00002e41;
power_data[313] = 32'h00002e41;
power_data[314] = 32'h00002e41;
power_data[315] = 32'h00002e41;
power_data[316] = 32'h00002e41;
power_data[317] = 32'h00002e41;
power_data[318] = 32'h00002e41;
power_data[319] = 32'h00002e41;
power_data[320] = 32'h00002e41;
power_data[321] = 32'h00002e41;
power_data[322] = 32'h00002e41;
power_data[323] = 32'h00002e41;
power_data[324] = 32'h00002e41;
power_data[325] = 32'h00002e41;
power_data[326] = 32'h00002e41;
power_data[327] = 32'h00002e41;
power_data[328] = 32'h00002e41;
power_data[329] = 32'h00002e41;
power_data[330] = 32'h00002e41;
power_data[331] = 32'h00002e41;
power_data[332] = 32'h00002e41;
power_data[333] = 32'h00002e41;
power_data[334] = 32'h00002e41;
power_data[335] = 32'h00002e41;
power_data[336] = 32'h00002e41;
power_data[337] = 32'h00002e41;
power_data[338] = 32'h00002e41;
power_data[339] = 32'h00002e41;
power_data[340] = 32'h00002e41;
power_data[341] = 32'h00002e41;
power_data[342] = 32'h00002e41;
power_data[343] = 32'h00002e41;
power_data[344] = 32'h00002e41;
power_data[345] = 32'h00002e41;
power_data[346] = 32'h00002e41;
power_data[347] = 32'h00002e41;
power_data[348] = 32'h00002e41;
power_data[349] = 32'h00002e41;
power_data[350] = 32'h00002e41;
power_data[351] = 32'h00002e41;
power_data[352] = 32'h00002e41;
power_data[353] = 32'h00002e41;
power_data[354] = 32'h000009ab;
power_data[355] = 32'h00000086;
power_data[356] = 32'h00000086;
power_data[357] = 32'h00000086;
power_data[358] = 32'h00000086;
power_data[359] = 32'h00000086;
power_data[360] = 32'h00000086;
power_data[361] = 32'h00000086;
power_data[362] = 32'h00000086;
power_data[363] = 32'h00000086;
power_data[364] = 32'h00000086;
power_data[365] = 32'h00000086;
power_data[366] = 32'h00000086;
power_data[367] = 32'h00000086;
power_data[368] = 32'h00000086;
power_data[369] = 32'h00000086;
power_data[370] = 32'h00000086;
power_data[371] = 32'h00000086;
power_data[372] = 32'h00000086;
power_data[373] = 32'h00000086;
power_data[374] = 32'h00000086;
power_data[375] = 32'h00000086;
power_data[376] = 32'h00000086;
power_data[377] = 32'h00000086;
power_data[378] = 32'h00000086;
power_data[379] = 32'h00000086;
power_data[380] = 32'h00000086;
power_data[381] = 32'h00000086;
power_data[382] = 32'h00000086;
power_data[383] = 32'h00000086;
power_data[384] = 32'h00000086;
power_data[385] = 32'h00000086;
power_data[386] = 32'h00000086;
power_data[387] = 32'h00000086;
power_data[388] = 32'h00000086;
power_data[389] = 32'h00000086;
power_data[390] = 32'h00000086;
power_data[391] = 32'h00000086;
power_data[392] = 32'h00000086;
power_data[393] = 32'h00000086;
power_data[394] = 32'h00000086;
power_data[395] = 32'h00000086;
power_data[396] = 32'h00000086;
power_data[397] = 32'h00000086;
power_data[398] = 32'h00000086;
power_data[399] = 32'h00000086;
power_data[400] = 32'h00000086;
power_data[401] = 32'h00000086;
power_data[402] = 32'h00000086;
power_data[403] = 32'h00000086;
power_data[404] = 32'h00000086;
power_data[405] = 32'h00000086;
power_data[406] = 32'h00000086;
power_data[407] = 32'h00000086;
power_data[408] = 32'h00000086;
power_data[409] = 32'h00000086;
power_data[410] = 32'h00000086;
power_data[411] = 32'h00000086;
power_data[412] = 32'h00000086;
power_data[413] = 32'h00000086;
power_data[414] = 32'h00000086;
power_data[415] = 32'h00000086;
power_data[416] = 32'h00000086;
power_data[417] = 32'h00000086;
power_data[418] = 32'h00000086;
power_data[419] = 32'h00000086;
power_data[420] = 32'h00000086;
power_data[421] = 32'h00000086;
power_data[422] = 32'h00000086;
power_data[423] = 32'h00000086;
power_data[424] = 32'h00000086;
power_data[425] = 32'h00000086;
power_data[426] = 32'h00000086;
power_data[427] = 32'h00000086;
power_data[428] = 32'h00000086;
power_data[429] = 32'h00000086;
power_data[430] = 32'h00000086;
power_data[431] = 32'h00000086;
power_data[432] = 32'h00000086;
power_data[433] = 32'h00000086;
power_data[434] = 32'h00000086;
power_data[435] = 32'h00000086;
power_data[436] = 32'h00000086;
power_data[437] = 32'h00000086;
power_data[438] = 32'h00000086;
power_data[439] = 32'h00000086;
power_data[440] = 32'h00000086;
power_data[441] = 32'h00000086;
power_data[442] = 32'h00000086;
power_data[443] = 32'h00000086;
power_data[444] = 32'h00000086;
power_data[445] = 32'h00000086;
power_data[446] = 32'h00000086;
power_data[447] = 32'h00000086;
power_data[448] = 32'h00000086;
power_data[449] = 32'h00000086;
power_data[450] = 32'h00000086;
power_data[451] = 32'h00000086;
power_data[452] = 32'h00000086;
power_data[453] = 32'h00000086;
power_data[454] = 32'h00000086;
power_data[455] = 32'h00000086;
power_data[456] = 32'h00000086;
power_data[457] = 32'h00000086;
power_data[458] = 32'h00000086;
power_data[459] = 32'h00000086;
power_data[460] = 32'h00000086;
power_data[461] = 32'h00000086;
power_data[462] = 32'h00000086;
power_data[463] = 32'h00000086;
power_data[464] = 32'h00000086;
power_data[465] = 32'h00000086;
power_data[466] = 32'h00000086;
power_data[467] = 32'h00000086;
power_data[468] = 32'h00000086;
power_data[469] = 32'h00000086;
power_data[470] = 32'h00000086;
power_data[471] = 32'h00000086;
power_data[472] = 32'h00000086;
power_data[473] = 32'h00000086;
power_data[474] = 32'h00000086;
power_data[475] = 32'h00000086;
power_data[476] = 32'h00000086;
power_data[477] = 32'h00000086;
power_data[478] = 32'h00000086;
power_data[479] = 32'h00000086;
power_data[480] = 32'h00000086;
power_data[481] = 32'h00000086;
power_data[482] = 32'h00000086;
power_data[483] = 32'h00000086;
power_data[484] = 32'h00000086;
power_data[485] = 32'h00000086;
power_data[486] = 32'h00000086;
power_data[487] = 32'h00000086;
power_data[488] = 32'h00000086;
power_data[489] = 32'h00000086;
power_data[490] = 32'h00000086;
power_data[491] = 32'h00000086;
power_data[492] = 32'h00000086;
power_data[493] = 32'h00000086;
power_data[494] = 32'h00000086;
power_data[495] = 32'h00000086;
power_data[496] = 32'h00000086;
power_data[497] = 32'h00000086;
power_data[498] = 32'h00000086;
power_data[499] = 32'h00000086;
power_data[500] = 32'h00000086;
power_data[501] = 32'h00000086;
power_data[502] = 32'h00000086;
power_data[503] = 32'h00000086;
power_data[504] = 32'h00000086;
power_data[505] = 32'h00000086;
power_data[506] = 32'h00000086;
power_data[507] = 32'h00000086;
power_data[508] = 32'h00000086;
power_data[509] = 32'h00000086;
power_data[510] = 32'h00000086;
power_data[511] = 32'h00000086;
power_data[512] = 32'h00000086;
power_data[513] = 32'h00000086;
power_data[514] = 32'h00000086;
power_data[515] = 32'h00000086;
power_data[516] = 32'h00000086;
power_data[517] = 32'h00000086;
power_data[518] = 32'h00000086;
power_data[519] = 32'h00000086;
power_data[520] = 32'h00000086;
power_data[521] = 32'h00000086;
power_data[522] = 32'h00000086;
power_data[523] = 32'h00000086;
power_data[524] = 32'h00000086;
power_data[525] = 32'h00000086;
power_data[526] = 32'h00000086;
power_data[527] = 32'h00000086;
power_data[528] = 32'h00000086;
power_data[529] = 32'h00000086;
power_data[530] = 32'h00000086;
power_data[531] = 32'h00000086;
power_data[532] = 32'h00000086;
power_data[533] = 32'h00000086;
power_data[534] = 32'h00000086;
power_data[535] = 32'h00000086;
power_data[536] = 32'h00000086;
power_data[537] = 32'h00000086;
power_data[538] = 32'h00000086;
power_data[539] = 32'h00000086;
power_data[540] = 32'h00000086;
power_data[541] = 32'h00000086;
power_data[542] = 32'h00000086;
power_data[543] = 32'h00000086;
power_data[544] = 32'h00000086;
power_data[545] = 32'h00000086;
power_data[546] = 32'h00000086;
power_data[547] = 32'h00000086;
power_data[548] = 32'h00000086;
power_data[549] = 32'h00000086;
power_data[550] = 32'h00000086;
power_data[551] = 32'h00000086;
power_data[552] = 32'h00000086;
power_data[553] = 32'h00000086;
power_data[554] = 32'h00000086;
power_data[555] = 32'h00000086;
power_data[556] = 32'h00000086;
power_data[557] = 32'h00000086;
power_data[558] = 32'h00000086;
power_data[559] = 32'h00000086;
power_data[560] = 32'h00000086;
power_data[561] = 32'h00000086;
power_data[562] = 32'h00000086;
power_data[563] = 32'h00000086;
power_data[564] = 32'h00000086;
power_data[565] = 32'h00000086;
power_data[566] = 32'h00000086;
power_data[567] = 32'h00000086;
power_data[568] = 32'h00000086;
power_data[569] = 32'h00000086;
power_data[570] = 32'h00000086;
power_data[571] = 32'h00000086;
power_data[572] = 32'h00000086;
power_data[573] = 32'h00000086;
power_data[574] = 32'h00000086;
power_data[575] = 32'h00000086;
power_data[576] = 32'h00000086;
power_data[577] = 32'h00000086;
power_data[578] = 32'h00000086;
power_data[579] = 32'h00000086;
power_data[580] = 32'h00000086;
power_data[581] = 32'h00000086;
power_data[582] = 32'h00000086;
power_data[583] = 32'h00000086;
power_data[584] = 32'h00000086;
power_data[585] = 32'h00000086;
power_data[586] = 32'h00000086;
power_data[587] = 32'h00000086;
power_data[588] = 32'h00000086;
power_data[589] = 32'h00000086;
power_data[590] = 32'h00000086;
power_data[591] = 32'h00000086;
power_data[592] = 32'h00000086;
power_data[593] = 32'h00000086;
power_data[594] = 32'h00000086;
power_data[595] = 32'h00000086;
power_data[596] = 32'h00000086;
power_data[597] = 32'h00000086;
power_data[598] = 32'h00000086;
power_data[599] = 32'h00000086;
power_data[600] = 32'h00000086;
power_data[601] = 32'h00000086;
power_data[602] = 32'h00000086;
power_data[603] = 32'h00000086;
power_data[604] = 32'h00000086;
power_data[605] = 32'h00000086;
power_data[606] = 32'h00000086;
power_data[607] = 32'h00000086;
power_data[608] = 32'h00000086;
power_data[609] = 32'h00000086;
power_data[610] = 32'h00000086;
power_data[611] = 32'h00000086;
power_data[612] = 32'h00000086;
power_data[613] = 32'h00000086;
power_data[614] = 32'h00000086;
power_data[615] = 32'h00000086;
power_data[616] = 32'h00000086;
power_data[617] = 32'h00000086;
power_data[618] = 32'h00000086;
power_data[619] = 32'h00000086;
power_data[620] = 32'h00000086;
power_data[621] = 32'h00000086;
power_data[622] = 32'h00000086;
power_data[623] = 32'h00000086;
power_data[624] = 32'h00000086;
power_data[625] = 32'h00000086;
power_data[626] = 32'h00000086;
power_data[627] = 32'h00000086;
power_data[628] = 32'h00000086;
power_data[629] = 32'h00000086;
power_data[630] = 32'h00000086;
power_data[631] = 32'h00000086;
power_data[632] = 32'h00000086;
power_data[633] = 32'h00000086;
power_data[634] = 32'h00000086;
power_data[635] = 32'h00000086;
power_data[636] = 32'h00000086;
power_data[637] = 32'h00000086;
power_data[638] = 32'h00000086;
power_data[639] = 32'h00000086;
power_data[640] = 32'h00000086;
power_data[641] = 32'h00000086;
power_data[642] = 32'h00000086;
power_data[643] = 32'h00000086;
power_data[644] = 32'h00000086;
power_data[645] = 32'h00000086;
power_data[646] = 32'h00000086;
power_data[647] = 32'h00000086;
power_data[648] = 32'h00000086;
power_data[649] = 32'h00000086;
power_data[650] = 32'h00000086;
power_data[651] = 32'h00000086;
power_data[652] = 32'h00000086;
power_data[653] = 32'h00000086;
power_data[654] = 32'h00000086;
power_data[655] = 32'h00000086;
power_data[656] = 32'h00000086;
power_data[657] = 32'h00000086;
power_data[658] = 32'h00000086;
power_data[659] = 32'h00000086;
power_data[660] = 32'h00000086;
power_data[661] = 32'h00000086;
power_data[662] = 32'h00000086;
power_data[663] = 32'h00000086;
power_data[664] = 32'h00000086;
power_data[665] = 32'h00000086;
power_data[666] = 32'h00000086;
power_data[667] = 32'h00000082;
power_data[668] = 32'h00000069;
power_data[669] = 32'h00000069;
power_data[670] = 32'h00000069;
power_data[671] = 32'h00000069;
power_data[672] = 32'h00000069;
power_data[673] = 32'h00000069;
power_data[674] = 32'h00000069;
power_data[675] = 32'h00000069;
power_data[676] = 32'h00000069;
power_data[677] = 32'h00000069;
power_data[678] = 32'h00000069;
power_data[679] = 32'h00000069;
power_data[680] = 32'h00000069;
power_data[681] = 32'h00000069;
power_data[682] = 32'h00000069;
power_data[683] = 32'h00000069;
power_data[684] = 32'h00000069;
power_data[685] = 32'h00000069;
power_data[686] = 32'h00000069;
power_data[687] = 32'h00000069;
power_data[688] = 32'h00000069;
power_data[689] = 32'h00000069;
power_data[690] = 32'h00000069;
power_data[691] = 32'h00000069;
power_data[692] = 32'h00000069;
power_data[693] = 32'h00000069;
power_data[694] = 32'h00000069;
power_data[695] = 32'h00000069;
power_data[696] = 32'h00000069;
power_data[697] = 32'h00000069;
power_data[698] = 32'h00000069;
power_data[699] = 32'h00000069;
power_data[700] = 32'h00000069;
power_data[701] = 32'h00000069;
power_data[702] = 32'h00000069;
power_data[703] = 32'h00000069;
power_data[704] = 32'h00000069;
power_data[705] = 32'h00000069;
power_data[706] = 32'h00000069;
power_data[707] = 32'h00000069;
power_data[708] = 32'h00000069;
power_data[709] = 32'h00000069;
power_data[710] = 32'h00000069;
power_data[711] = 32'h00000069;
power_data[712] = 32'h00000069;
power_data[713] = 32'h00000069;
power_data[714] = 32'h00000069;
power_data[715] = 32'h00000069;
power_data[716] = 32'h00000069;
power_data[717] = 32'h00000069;
power_data[718] = 32'h00000069;
power_data[719] = 32'h00000069;
power_data[720] = 32'h00000069;
power_data[721] = 32'h00000069;
power_data[722] = 32'h00000069;
power_data[723] = 32'h00000069;
power_data[724] = 32'h00000069;
power_data[725] = 32'h00000069;
power_data[726] = 32'h00000069;
power_data[727] = 32'h00000069;
power_data[728] = 32'h00000069;
power_data[729] = 32'h00000069;
power_data[730] = 32'h00000069;
power_data[731] = 32'h00000069;
power_data[732] = 32'h00000069;
power_data[733] = 32'h00000069;
power_data[734] = 32'h00000069;
power_data[735] = 32'h00000069;
power_data[736] = 32'h00000069;
power_data[737] = 32'h00000069;
power_data[738] = 32'h0000077d;
power_data[739] = 32'h00000942;
power_data[740] = 32'h00000942;
power_data[741] = 32'h00000942;
power_data[742] = 32'h00000942;
power_data[743] = 32'h00000942;
power_data[744] = 32'h00000942;
power_data[745] = 32'h00000942;
power_data[746] = 32'h00000942;
power_data[747] = 32'h00000942;
power_data[748] = 32'h00000942;
power_data[749] = 32'h00000942;
power_data[750] = 32'h00000942;
power_data[751] = 32'h00000942;
power_data[752] = 32'h00000942;
power_data[753] = 32'h00000942;
power_data[754] = 32'h00000942;
power_data[755] = 32'h00000942;
power_data[756] = 32'h00000942;
power_data[757] = 32'h00000942;
power_data[758] = 32'h00000942;
power_data[759] = 32'h00000942;
power_data[760] = 32'h00000942;
power_data[761] = 32'h00000942;
power_data[762] = 32'h00000942;
power_data[763] = 32'h00000942;
power_data[764] = 32'h00000942;
power_data[765] = 32'h00000942;
power_data[766] = 32'h00000942;
power_data[767] = 32'h00000232;
power_data[768] = 32'h00000232;
power_data[769] = 32'h00000232;
power_data[770] = 32'h00000232;
power_data[771] = 32'h00000232;
power_data[772] = 32'h00000232;
power_data[773] = 32'h00000232;
power_data[774] = 32'h00000232;
power_data[775] = 32'h00000232;
power_data[776] = 32'h00000232;
power_data[777] = 32'h00000232;
power_data[778] = 32'h00000232;
power_data[779] = 32'h00000232;
power_data[780] = 32'h00000232;
power_data[781] = 32'h00000232;
power_data[782] = 32'h00000232;
power_data[783] = 32'h00000232;
power_data[784] = 32'h00000232;
power_data[785] = 32'h00000232;
power_data[786] = 32'h00000232;
power_data[787] = 32'h00000232;
power_data[788] = 32'h00000232;
power_data[789] = 32'h00000232;
power_data[790] = 32'h00000232;
power_data[791] = 32'h00000232;
power_data[792] = 32'h00000232;
power_data[793] = 32'h00000232;
power_data[794] = 32'h00000232;
power_data[795] = 32'h00000232;
power_data[796] = 32'h00000232;
power_data[797] = 32'h00000232;
power_data[798] = 32'h00000232;
power_data[799] = 32'h00000232;
power_data[800] = 32'h00000232;
power_data[801] = 32'h00000232;
power_data[802] = 32'h00000232;
power_data[803] = 32'h00000232;
power_data[804] = 32'h00000232;
power_data[805] = 32'h00000232;
power_data[806] = 32'h00000232;
power_data[807] = 32'h00000232;
power_data[808] = 32'h000013d3;
power_data[809] = 32'h00002e41;
power_data[810] = 32'h00002e41;
power_data[811] = 32'h00002e41;
power_data[812] = 32'h00002e41;
power_data[813] = 32'h00002e41;
power_data[814] = 32'h00002e41;
power_data[815] = 32'h00002e41;
power_data[816] = 32'h00002e41;
power_data[817] = 32'h00002e41;
power_data[818] = 32'h00002e41;
power_data[819] = 32'h00002e41;
power_data[820] = 32'h00002e41;
power_data[821] = 32'h00002e41;
power_data[822] = 32'h00002e41;
power_data[823] = 32'h00002e41;
power_data[824] = 32'h00002e41;
power_data[825] = 32'h00002e41;
power_data[826] = 32'h00002e41;
power_data[827] = 32'h00002e41;
power_data[828] = 32'h00002e41;
power_data[829] = 32'h00002e41;
power_data[830] = 32'h00002e41;
power_data[831] = 32'h00002e41;
power_data[832] = 32'h00002e41;
power_data[833] = 32'h00002e41;
power_data[834] = 32'h00002e41;
power_data[835] = 32'h00002e41;
power_data[836] = 32'h00002e41;
power_data[837] = 32'h00002e41;
power_data[838] = 32'h00002e41;
power_data[839] = 32'h00002e41;
power_data[840] = 32'h00002e41;
power_data[841] = 32'h00002e41;
power_data[842] = 32'h00002e41;
power_data[843] = 32'h00002e41;
power_data[844] = 32'h00002e41;
power_data[845] = 32'h00002e41;
power_data[846] = 32'h00002e41;
power_data[847] = 32'h00002e41;
power_data[848] = 32'h00002e41;
power_data[849] = 32'h00002e41;
power_data[850] = 32'h00002e41;
power_data[851] = 32'h00002e41;
power_data[852] = 32'h00002e41;
power_data[853] = 32'h00002e41;
power_data[854] = 32'h00002e41;
power_data[855] = 32'h00002e41;
power_data[856] = 32'h00002e41;
power_data[857] = 32'h00002e41;
power_data[858] = 32'h00002e41;
power_data[859] = 32'h00002e41;
power_data[860] = 32'h00002e41;
power_data[861] = 32'h00002e41;
power_data[862] = 32'h00002e41;
power_data[863] = 32'h00002e41;
power_data[864] = 32'h00002e41;
power_data[865] = 32'h00002e41;
power_data[866] = 32'h000009ab;
power_data[867] = 32'h00000086;
power_data[868] = 32'h00000086;
power_data[869] = 32'h00000086;
power_data[870] = 32'h00000086;
power_data[871] = 32'h00000086;
power_data[872] = 32'h00000086;
power_data[873] = 32'h00000086;
power_data[874] = 32'h00000086;
power_data[875] = 32'h00000086;
power_data[876] = 32'h00000086;
power_data[877] = 32'h00000086;
power_data[878] = 32'h00000086;
power_data[879] = 32'h00000086;
power_data[880] = 32'h00000086;
power_data[881] = 32'h00000086;
power_data[882] = 32'h00000086;
power_data[883] = 32'h00000086;
power_data[884] = 32'h00000086;
power_data[885] = 32'h00000086;
power_data[886] = 32'h00000086;
power_data[887] = 32'h00000086;
power_data[888] = 32'h00000086;
power_data[889] = 32'h00000086;
power_data[890] = 32'h00000086;
power_data[891] = 32'h00000086;
power_data[892] = 32'h00000086;
power_data[893] = 32'h00000086;
power_data[894] = 32'h00000086;
power_data[895] = 32'h00000086;
power_data[896] = 32'h00000086;
power_data[897] = 32'h00000086;
power_data[898] = 32'h00000086;
power_data[899] = 32'h00000086;
power_data[900] = 32'h00000086;
power_data[901] = 32'h00000086;
power_data[902] = 32'h00000086;
power_data[903] = 32'h00000086;
power_data[904] = 32'h00000086;
power_data[905] = 32'h00000086;
power_data[906] = 32'h00000086;
power_data[907] = 32'h00000086;
power_data[908] = 32'h00000086;
power_data[909] = 32'h00000086;
power_data[910] = 32'h00000086;
power_data[911] = 32'h00000086;
power_data[912] = 32'h00000086;
power_data[913] = 32'h00000086;
power_data[914] = 32'h00000086;
power_data[915] = 32'h00000086;
power_data[916] = 32'h00000086;
power_data[917] = 32'h00000086;
power_data[918] = 32'h00000086;
power_data[919] = 32'h00000086;
power_data[920] = 32'h00000086;
power_data[921] = 32'h00000086;
power_data[922] = 32'h00000086;
power_data[923] = 32'h00000086;
power_data[924] = 32'h00000086;
power_data[925] = 32'h00000086;
power_data[926] = 32'h00000086;
power_data[927] = 32'h00000086;
power_data[928] = 32'h00000086;
power_data[929] = 32'h00000086;
power_data[930] = 32'h00000086;
power_data[931] = 32'h00000086;
power_data[932] = 32'h00000086;
power_data[933] = 32'h00000086;
power_data[934] = 32'h00000086;
power_data[935] = 32'h00000086;
power_data[936] = 32'h00000086;
power_data[937] = 32'h00000086;
power_data[938] = 32'h00000086;
power_data[939] = 32'h00000086;
power_data[940] = 32'h00000086;
power_data[941] = 32'h00000086;
power_data[942] = 32'h00000086;
power_data[943] = 32'h00000086;
power_data[944] = 32'h00000086;
power_data[945] = 32'h00000086;
power_data[946] = 32'h00000086;
power_data[947] = 32'h00000086;
power_data[948] = 32'h00000086;
power_data[949] = 32'h00000086;
power_data[950] = 32'h00000086;
power_data[951] = 32'h00000086;
power_data[952] = 32'h00000086;
power_data[953] = 32'h00000086;
power_data[954] = 32'h00000086;
power_data[955] = 32'h00000086;
power_data[956] = 32'h00000086;
power_data[957] = 32'h00000086;
power_data[958] = 32'h00000086;
power_data[959] = 32'h00000086;
power_data[960] = 32'h00000086;
power_data[961] = 32'h00000086;
power_data[962] = 32'h00000086;
power_data[963] = 32'h00000086;
power_data[964] = 32'h00000086;
power_data[965] = 32'h00000086;
power_data[966] = 32'h00000086;
power_data[967] = 32'h00000086;
power_data[968] = 32'h00000086;
power_data[969] = 32'h00000086;
power_data[970] = 32'h00000086;
power_data[971] = 32'h00000086;
power_data[972] = 32'h00000086;
power_data[973] = 32'h00000086;
power_data[974] = 32'h00000086;
power_data[975] = 32'h00000086;
power_data[976] = 32'h00000086;
power_data[977] = 32'h00000086;
power_data[978] = 32'h00000086;
power_data[979] = 32'h00000086;
power_data[980] = 32'h00000086;
power_data[981] = 32'h00000086;
power_data[982] = 32'h00000086;
power_data[983] = 32'h00000086;
power_data[984] = 32'h00000086;
power_data[985] = 32'h00000086;
power_data[986] = 32'h00000086;
power_data[987] = 32'h00000086;
power_data[988] = 32'h00000086;
power_data[989] = 32'h00000086;
power_data[990] = 32'h00000086;
power_data[991] = 32'h00000086;
power_data[992] = 32'h00000086;
power_data[993] = 32'h00000086;
power_data[994] = 32'h00000086;
power_data[995] = 32'h00000086;
power_data[996] = 32'h00000086;
power_data[997] = 32'h00000086;
power_data[998] = 32'h00000086;
power_data[999] = 32'h00000086;
power_data[1000] = 32'h00000086;
power_data[1001] = 32'h00000086;
power_data[1002] = 32'h00000086;
power_data[1003] = 32'h00000086;
power_data[1004] = 32'h00000086;
power_data[1005] = 32'h00000086;
power_data[1006] = 32'h00000086;
power_data[1007] = 32'h00000086;
power_data[1008] = 32'h00000086;
power_data[1009] = 32'h00000086;
power_data[1010] = 32'h00000086;
power_data[1011] = 32'h00000086;
power_data[1012] = 32'h00000086;
power_data[1013] = 32'h00000086;
power_data[1014] = 32'h00000086;
power_data[1015] = 32'h00000086;
power_data[1016] = 32'h00000086;
power_data[1017] = 32'h00000086;
power_data[1018] = 32'h00000086;
power_data[1019] = 32'h00000086;
power_data[1020] = 32'h00000086;
power_data[1021] = 32'h00000086;
power_data[1022] = 32'h00000086;
power_data[1023] = 32'h00000086;
power_data[1024] = 32'h00000086;
power_data[1025] = 32'h00000086;
power_data[1026] = 32'h00000086;
power_data[1027] = 32'h00000086;
power_data[1028] = 32'h00000086;
power_data[1029] = 32'h00000086;
power_data[1030] = 32'h00000086;
power_data[1031] = 32'h00000086;
power_data[1032] = 32'h00000086;
power_data[1033] = 32'h00000086;
power_data[1034] = 32'h00000086;
power_data[1035] = 32'h00000086;
power_data[1036] = 32'h00000086;
power_data[1037] = 32'h00000086;
power_data[1038] = 32'h00000086;
power_data[1039] = 32'h00000086;
power_data[1040] = 32'h00000086;
power_data[1041] = 32'h00000086;
power_data[1042] = 32'h00000086;
power_data[1043] = 32'h00000086;
power_data[1044] = 32'h00000086;
power_data[1045] = 32'h00000086;
power_data[1046] = 32'h00000086;
power_data[1047] = 32'h00000086;
power_data[1048] = 32'h00000086;
power_data[1049] = 32'h00000086;
power_data[1050] = 32'h00000086;
power_data[1051] = 32'h00000086;
power_data[1052] = 32'h00000086;
power_data[1053] = 32'h00000086;
power_data[1054] = 32'h00000086;
power_data[1055] = 32'h00000086;
power_data[1056] = 32'h00000086;
power_data[1057] = 32'h00000086;
power_data[1058] = 32'h00000086;
power_data[1059] = 32'h00000086;
power_data[1060] = 32'h00000086;
power_data[1061] = 32'h00000086;
power_data[1062] = 32'h00000086;
power_data[1063] = 32'h00000086;
power_data[1064] = 32'h00000086;
power_data[1065] = 32'h00000086;
power_data[1066] = 32'h00000086;
power_data[1067] = 32'h00000086;
power_data[1068] = 32'h00000086;
power_data[1069] = 32'h00000086;
power_data[1070] = 32'h00000086;
power_data[1071] = 32'h00000086;
power_data[1072] = 32'h00000086;
power_data[1073] = 32'h00000086;
power_data[1074] = 32'h00000086;
power_data[1075] = 32'h00000086;
power_data[1076] = 32'h00000086;
power_data[1077] = 32'h00000086;
power_data[1078] = 32'h00000086;
power_data[1079] = 32'h00000086;
power_data[1080] = 32'h00000086;
power_data[1081] = 32'h00000086;
power_data[1082] = 32'h00000086;
power_data[1083] = 32'h00000086;
power_data[1084] = 32'h00000086;
power_data[1085] = 32'h00000086;
power_data[1086] = 32'h00000086;
power_data[1087] = 32'h00000086;
power_data[1088] = 32'h00000086;
power_data[1089] = 32'h00000086;
power_data[1090] = 32'h00000086;
power_data[1091] = 32'h00000086;
power_data[1092] = 32'h00000086;
power_data[1093] = 32'h00000086;
power_data[1094] = 32'h00000086;
power_data[1095] = 32'h00000086;
power_data[1096] = 32'h00000086;
power_data[1097] = 32'h00000086;
power_data[1098] = 32'h00000086;
power_data[1099] = 32'h00000086;
power_data[1100] = 32'h00000086;
power_data[1101] = 32'h00000086;
power_data[1102] = 32'h00000086;
power_data[1103] = 32'h00000086;
power_data[1104] = 32'h00000086;
power_data[1105] = 32'h00000086;
power_data[1106] = 32'h00000086;
power_data[1107] = 32'h00000086;
power_data[1108] = 32'h00000086;
power_data[1109] = 32'h00000086;
power_data[1110] = 32'h00000086;
power_data[1111] = 32'h00000086;
power_data[1112] = 32'h00000086;
power_data[1113] = 32'h00000086;
power_data[1114] = 32'h00000086;
power_data[1115] = 32'h00000086;
power_data[1116] = 32'h00000086;
power_data[1117] = 32'h00000086;
power_data[1118] = 32'h00000086;
power_data[1119] = 32'h00000086;
power_data[1120] = 32'h00000086;
power_data[1121] = 32'h00000086;
power_data[1122] = 32'h00000086;
power_data[1123] = 32'h00000086;
power_data[1124] = 32'h00000086;
power_data[1125] = 32'h00000086;
power_data[1126] = 32'h00000086;
power_data[1127] = 32'h00000086;
power_data[1128] = 32'h00000086;
power_data[1129] = 32'h00000086;
power_data[1130] = 32'h00000086;
power_data[1131] = 32'h00000086;
power_data[1132] = 32'h00000086;
power_data[1133] = 32'h00000086;
power_data[1134] = 32'h00000086;
power_data[1135] = 32'h00000086;
power_data[1136] = 32'h00000086;
power_data[1137] = 32'h00000086;
power_data[1138] = 32'h00000086;
power_data[1139] = 32'h00000086;
power_data[1140] = 32'h00000086;
power_data[1141] = 32'h00000086;
power_data[1142] = 32'h00000086;
power_data[1143] = 32'h00000086;
power_data[1144] = 32'h00000086;
power_data[1145] = 32'h00000086;
power_data[1146] = 32'h00000086;
power_data[1147] = 32'h00000086;
power_data[1148] = 32'h00000086;
power_data[1149] = 32'h00000086;
power_data[1150] = 32'h00000086;
power_data[1151] = 32'h00000086;
power_data[1152] = 32'h00000086;
power_data[1153] = 32'h00000086;
power_data[1154] = 32'h00000086;
power_data[1155] = 32'h00000086;
power_data[1156] = 32'h00000086;
power_data[1157] = 32'h00000086;
power_data[1158] = 32'h00000086;
power_data[1159] = 32'h00000086;
power_data[1160] = 32'h00000086;
power_data[1161] = 32'h00000086;
power_data[1162] = 32'h00000086;
power_data[1163] = 32'h00000086;
power_data[1164] = 32'h00000086;
power_data[1165] = 32'h00000086;
power_data[1166] = 32'h00000086;
power_data[1167] = 32'h00000086;
power_data[1168] = 32'h00000086;
power_data[1169] = 32'h00000086;
power_data[1170] = 32'h00000086;
power_data[1171] = 32'h00000086;
power_data[1172] = 32'h00000086;
power_data[1173] = 32'h00000086;
power_data[1174] = 32'h00000086;
power_data[1175] = 32'h00000086;
power_data[1176] = 32'h00000086;
power_data[1177] = 32'h00000086;
power_data[1178] = 32'h00000086;
power_data[1179] = 32'h00000082;
power_data[1180] = 32'h00000069;
power_data[1181] = 32'h00000069;
power_data[1182] = 32'h00000069;
power_data[1183] = 32'h00000069;
power_data[1184] = 32'h00000069;
power_data[1185] = 32'h00000069;
power_data[1186] = 32'h00000069;
power_data[1187] = 32'h00000069;
power_data[1188] = 32'h00000069;
power_data[1189] = 32'h00000069;
power_data[1190] = 32'h00000069;
power_data[1191] = 32'h00000069;
power_data[1192] = 32'h00000069;
power_data[1193] = 32'h00000069;
power_data[1194] = 32'h00000069;
power_data[1195] = 32'h00000069;
power_data[1196] = 32'h00000069;
power_data[1197] = 32'h00000069;
power_data[1198] = 32'h00000069;
power_data[1199] = 32'h00000069;
power_data[1200] = 32'h00000069;
power_data[1201] = 32'h00000069;
power_data[1202] = 32'h00000069;
power_data[1203] = 32'h00000069;
power_data[1204] = 32'h00000069;
power_data[1205] = 32'h00000069;
power_data[1206] = 32'h00000069;
power_data[1207] = 32'h00000069;
power_data[1208] = 32'h00000069;
power_data[1209] = 32'h00000069;
power_data[1210] = 32'h00000069;
power_data[1211] = 32'h00000069;
power_data[1212] = 32'h00000069;
power_data[1213] = 32'h00000069;
power_data[1214] = 32'h00000069;
power_data[1215] = 32'h00000069;
power_data[1216] = 32'h00000069;
power_data[1217] = 32'h00000069;
power_data[1218] = 32'h00000069;
power_data[1219] = 32'h00000069;
power_data[1220] = 32'h00000069;
power_data[1221] = 32'h00000069;
power_data[1222] = 32'h00000069;
power_data[1223] = 32'h00000069;
power_data[1224] = 32'h00000069;
power_data[1225] = 32'h00000069;
power_data[1226] = 32'h00000069;
power_data[1227] = 32'h00000069;
power_data[1228] = 32'h00000069;
power_data[1229] = 32'h00000069;
power_data[1230] = 32'h00000069;
power_data[1231] = 32'h00000069;
power_data[1232] = 32'h00000069;
power_data[1233] = 32'h00000069;
power_data[1234] = 32'h00000069;
power_data[1235] = 32'h00000069;
power_data[1236] = 32'h00000069;
power_data[1237] = 32'h00000069;
power_data[1238] = 32'h00000069;
power_data[1239] = 32'h00000069;
power_data[1240] = 32'h00000069;
power_data[1241] = 32'h00000069;
power_data[1242] = 32'h00000069;
power_data[1243] = 32'h00000069;
power_data[1244] = 32'h00000069;
power_data[1245] = 32'h00000069;
power_data[1246] = 32'h00000069;
power_data[1247] = 32'h00000069;
power_data[1248] = 32'h00000069;
power_data[1249] = 32'h00000069;
power_data[1250] = 32'h0000077d;
power_data[1251] = 32'h00000942;
power_data[1252] = 32'h00000942;
power_data[1253] = 32'h00000942;
power_data[1254] = 32'h00000942;
power_data[1255] = 32'h00000942;
power_data[1256] = 32'h00000942;
power_data[1257] = 32'h00000942;
power_data[1258] = 32'h00000942;
power_data[1259] = 32'h00000942;
power_data[1260] = 32'h00000942;
power_data[1261] = 32'h00000942;
power_data[1262] = 32'h00000942;
power_data[1263] = 32'h00000942;
power_data[1264] = 32'h00000942;
power_data[1265] = 32'h00000942;
power_data[1266] = 32'h00000942;
power_data[1267] = 32'h00000942;
power_data[1268] = 32'h00000942;
power_data[1269] = 32'h00000942;
power_data[1270] = 32'h00000942;
power_data[1271] = 32'h00000942;
power_data[1272] = 32'h00000942;
power_data[1273] = 32'h00000942;
power_data[1274] = 32'h00000942;
power_data[1275] = 32'h00000942;
power_data[1276] = 32'h00000942;
power_data[1277] = 32'h00000942;
power_data[1278] = 32'h00000942;
power_data[1279] = 32'h00000232;
power_data[1280] = 32'h00000232;
power_data[1281] = 32'h00000232;
power_data[1282] = 32'h00000232;
power_data[1283] = 32'h00000232;
power_data[1284] = 32'h00000232;
power_data[1285] = 32'h00000232;
power_data[1286] = 32'h00000232;
power_data[1287] = 32'h00000232;
power_data[1288] = 32'h00000232;
power_data[1289] = 32'h00000232;
power_data[1290] = 32'h00000232;
power_data[1291] = 32'h00000232;
power_data[1292] = 32'h00000232;
power_data[1293] = 32'h00000232;
power_data[1294] = 32'h00000232;
power_data[1295] = 32'h00000232;
power_data[1296] = 32'h00000232;
power_data[1297] = 32'h00000232;
power_data[1298] = 32'h00000232;
power_data[1299] = 32'h00000232;
power_data[1300] = 32'h00000232;
power_data[1301] = 32'h00000232;
power_data[1302] = 32'h00000232;
power_data[1303] = 32'h00000232;
power_data[1304] = 32'h00000232;
power_data[1305] = 32'h00000232;
power_data[1306] = 32'h00000232;
power_data[1307] = 32'h00000232;
power_data[1308] = 32'h00000232;
power_data[1309] = 32'h00000232;
power_data[1310] = 32'h00000232;
power_data[1311] = 32'h00000232;
power_data[1312] = 32'h00000232;
power_data[1313] = 32'h00000232;
power_data[1314] = 32'h00000232;
power_data[1315] = 32'h00000232;
power_data[1316] = 32'h00000232;
power_data[1317] = 32'h00000232;
power_data[1318] = 32'h00000232;
power_data[1319] = 32'h00000232;
power_data[1320] = 32'h000013d3;
power_data[1321] = 32'h00002e41;
power_data[1322] = 32'h00002e41;
power_data[1323] = 32'h00002e41;
power_data[1324] = 32'h00002e41;
power_data[1325] = 32'h00002e41;
power_data[1326] = 32'h00002e41;
power_data[1327] = 32'h00002e41;
power_data[1328] = 32'h00002e41;
power_data[1329] = 32'h00002e41;
power_data[1330] = 32'h00002e41;
power_data[1331] = 32'h00002e41;
power_data[1332] = 32'h00002e41;
power_data[1333] = 32'h00002e41;
power_data[1334] = 32'h00002e41;
power_data[1335] = 32'h00002e41;
power_data[1336] = 32'h00002e41;
power_data[1337] = 32'h00002e41;
power_data[1338] = 32'h00002e41;
power_data[1339] = 32'h00002e41;
power_data[1340] = 32'h00002e41;
power_data[1341] = 32'h00002e41;
power_data[1342] = 32'h00002e41;
power_data[1343] = 32'h00002e41;
power_data[1344] = 32'h00002e41;
power_data[1345] = 32'h00002e41;
power_data[1346] = 32'h00002e41;
power_data[1347] = 32'h00002e41;
power_data[1348] = 32'h00002e41;
power_data[1349] = 32'h00002e41;
power_data[1350] = 32'h00002e41;
power_data[1351] = 32'h00002e41;
power_data[1352] = 32'h00002e41;
power_data[1353] = 32'h00002e41;
power_data[1354] = 32'h00002e41;
power_data[1355] = 32'h00002e41;
power_data[1356] = 32'h00002e41;
power_data[1357] = 32'h00002e41;
power_data[1358] = 32'h00002e41;
power_data[1359] = 32'h00002e41;
power_data[1360] = 32'h00002e41;
power_data[1361] = 32'h00002e41;
power_data[1362] = 32'h00002e41;
power_data[1363] = 32'h00002e41;
power_data[1364] = 32'h00002e41;
power_data[1365] = 32'h00002e41;
power_data[1366] = 32'h00002e41;
power_data[1367] = 32'h00002e41;
power_data[1368] = 32'h00002e41;
power_data[1369] = 32'h00002e41;
power_data[1370] = 32'h00002e41;
power_data[1371] = 32'h00002e41;
power_data[1372] = 32'h00002e41;
power_data[1373] = 32'h00002e41;
power_data[1374] = 32'h00002e41;
power_data[1375] = 32'h00002e41;
power_data[1376] = 32'h00002e41;
power_data[1377] = 32'h00002e41;
power_data[1378] = 32'h000009ab;
power_data[1379] = 32'h00000086;
power_data[1380] = 32'h00000086;
power_data[1381] = 32'h00000086;
power_data[1382] = 32'h00000086;
power_data[1383] = 32'h00000086;
power_data[1384] = 32'h00000086;
power_data[1385] = 32'h00000086;
power_data[1386] = 32'h00000086;
power_data[1387] = 32'h00000086;
power_data[1388] = 32'h00000086;
power_data[1389] = 32'h00000086;
power_data[1390] = 32'h00000086;
power_data[1391] = 32'h00000086;
power_data[1392] = 32'h00000086;
power_data[1393] = 32'h00000086;
power_data[1394] = 32'h00000086;
power_data[1395] = 32'h00000086;
power_data[1396] = 32'h00000086;
power_data[1397] = 32'h00000086;
power_data[1398] = 32'h00000086;
power_data[1399] = 32'h00000086;
power_data[1400] = 32'h00000086;
power_data[1401] = 32'h00000086;
power_data[1402] = 32'h00000086;
power_data[1403] = 32'h00000086;
power_data[1404] = 32'h00000086;
power_data[1405] = 32'h00000086;
power_data[1406] = 32'h00000086;
power_data[1407] = 32'h00000086;
power_data[1408] = 32'h00000086;
power_data[1409] = 32'h00000086;
power_data[1410] = 32'h00000086;
power_data[1411] = 32'h00000086;
power_data[1412] = 32'h00000086;
power_data[1413] = 32'h00000086;
power_data[1414] = 32'h00000086;
power_data[1415] = 32'h00000086;
power_data[1416] = 32'h00000086;
power_data[1417] = 32'h00000086;
power_data[1418] = 32'h00000086;
power_data[1419] = 32'h00000086;
power_data[1420] = 32'h00000086;
power_data[1421] = 32'h00000086;
power_data[1422] = 32'h00000086;
power_data[1423] = 32'h00000086;
power_data[1424] = 32'h00000086;
power_data[1425] = 32'h00000086;
power_data[1426] = 32'h00000086;
power_data[1427] = 32'h00000086;
power_data[1428] = 32'h00000086;
power_data[1429] = 32'h00000086;
power_data[1430] = 32'h00000086;
power_data[1431] = 32'h00000086;
power_data[1432] = 32'h00000086;
power_data[1433] = 32'h00000086;
power_data[1434] = 32'h00000086;
power_data[1435] = 32'h00000086;
power_data[1436] = 32'h00000086;
power_data[1437] = 32'h00000086;
power_data[1438] = 32'h00000086;
power_data[1439] = 32'h00000086;
power_data[1440] = 32'h00000086;
power_data[1441] = 32'h00000086;
power_data[1442] = 32'h00000086;
power_data[1443] = 32'h00000086;
power_data[1444] = 32'h00000086;
power_data[1445] = 32'h00000086;
power_data[1446] = 32'h00000086;
power_data[1447] = 32'h00000086;
power_data[1448] = 32'h00000086;
power_data[1449] = 32'h00000086;
power_data[1450] = 32'h00000086;
power_data[1451] = 32'h00000086;
power_data[1452] = 32'h00000086;
power_data[1453] = 32'h00000086;
power_data[1454] = 32'h00000086;
power_data[1455] = 32'h00000086;
power_data[1456] = 32'h00000086;
power_data[1457] = 32'h00000086;
power_data[1458] = 32'h00000086;
power_data[1459] = 32'h00000086;
power_data[1460] = 32'h00000086;
power_data[1461] = 32'h00000086;
power_data[1462] = 32'h00000086;
power_data[1463] = 32'h00000086;
power_data[1464] = 32'h00000086;
power_data[1465] = 32'h00000086;
power_data[1466] = 32'h00000086;
power_data[1467] = 32'h00000086;
power_data[1468] = 32'h00000086;
power_data[1469] = 32'h00000086;
power_data[1470] = 32'h00000086;
power_data[1471] = 32'h00000086;
power_data[1472] = 32'h00000086;
power_data[1473] = 32'h00000086;
power_data[1474] = 32'h00000086;
power_data[1475] = 32'h00000086;
power_data[1476] = 32'h00000086;
power_data[1477] = 32'h00000086;
power_data[1478] = 32'h00000086;
power_data[1479] = 32'h00000086;
power_data[1480] = 32'h00000086;
power_data[1481] = 32'h00000086;
power_data[1482] = 32'h00000086;
power_data[1483] = 32'h00000086;
power_data[1484] = 32'h00000086;
power_data[1485] = 32'h00000086;
power_data[1486] = 32'h00000086;
power_data[1487] = 32'h00000086;
power_data[1488] = 32'h00000086;
power_data[1489] = 32'h00000086;
power_data[1490] = 32'h00000086;
power_data[1491] = 32'h00000086;
power_data[1492] = 32'h00000086;
power_data[1493] = 32'h00000086;
power_data[1494] = 32'h00000086;
power_data[1495] = 32'h00000086;
power_data[1496] = 32'h00000086;
power_data[1497] = 32'h00000086;
power_data[1498] = 32'h00000086;
power_data[1499] = 32'h00000086;
power_data[1500] = 32'h00000086;
power_data[1501] = 32'h00000086;
power_data[1502] = 32'h00000086;
power_data[1503] = 32'h00000086;
power_data[1504] = 32'h00000086;
power_data[1505] = 32'h00000086;
power_data[1506] = 32'h00000086;
power_data[1507] = 32'h00000086;
power_data[1508] = 32'h00000086;
power_data[1509] = 32'h00000086;
power_data[1510] = 32'h00000086;
power_data[1511] = 32'h00000086;
power_data[1512] = 32'h00000086;
power_data[1513] = 32'h00000086;
power_data[1514] = 32'h00000086;
power_data[1515] = 32'h00000086;
power_data[1516] = 32'h00000086;
power_data[1517] = 32'h00000086;
power_data[1518] = 32'h00000086;
power_data[1519] = 32'h00000086;
power_data[1520] = 32'h00000086;
power_data[1521] = 32'h00000086;
power_data[1522] = 32'h00000086;
power_data[1523] = 32'h00000086;
power_data[1524] = 32'h00000086;
power_data[1525] = 32'h00000086;
power_data[1526] = 32'h00000086;
power_data[1527] = 32'h00000086;
power_data[1528] = 32'h00000086;
power_data[1529] = 32'h00000086;
power_data[1530] = 32'h00000086;
power_data[1531] = 32'h00000086;
power_data[1532] = 32'h00000086;
power_data[1533] = 32'h00000086;
power_data[1534] = 32'h00000086;
power_data[1535] = 32'h00000086;
power_data[1536] = 32'h00000086;
power_data[1537] = 32'h00000086;
power_data[1538] = 32'h00000086;
power_data[1539] = 32'h00000086;
power_data[1540] = 32'h00000086;
power_data[1541] = 32'h00000086;
power_data[1542] = 32'h00000086;
power_data[1543] = 32'h00000086;
power_data[1544] = 32'h00000086;
power_data[1545] = 32'h00000086;
power_data[1546] = 32'h00000086;
power_data[1547] = 32'h00000086;
power_data[1548] = 32'h00000086;
power_data[1549] = 32'h00000086;
power_data[1550] = 32'h00000086;
power_data[1551] = 32'h00000086;
power_data[1552] = 32'h00000086;
power_data[1553] = 32'h00000086;
power_data[1554] = 32'h00000086;
power_data[1555] = 32'h00000086;
power_data[1556] = 32'h00000086;
power_data[1557] = 32'h00000086;
power_data[1558] = 32'h00000086;
power_data[1559] = 32'h00000086;
power_data[1560] = 32'h00000086;
power_data[1561] = 32'h00000086;
power_data[1562] = 32'h00000086;
power_data[1563] = 32'h00000086;
power_data[1564] = 32'h00000086;
power_data[1565] = 32'h00000086;
power_data[1566] = 32'h00000086;
power_data[1567] = 32'h00000086;
power_data[1568] = 32'h00000086;
power_data[1569] = 32'h00000086;
power_data[1570] = 32'h00000086;
power_data[1571] = 32'h00000086;
power_data[1572] = 32'h00000086;
power_data[1573] = 32'h00000086;
power_data[1574] = 32'h00000086;
power_data[1575] = 32'h00000086;
power_data[1576] = 32'h00000086;
power_data[1577] = 32'h00000086;
power_data[1578] = 32'h00000086;
power_data[1579] = 32'h00000086;
power_data[1580] = 32'h00000086;
power_data[1581] = 32'h00000086;
power_data[1582] = 32'h00000086;
power_data[1583] = 32'h00000086;
power_data[1584] = 32'h00000086;
power_data[1585] = 32'h00000086;
power_data[1586] = 32'h00000086;
power_data[1587] = 32'h00000086;
power_data[1588] = 32'h00000086;
power_data[1589] = 32'h00000086;
power_data[1590] = 32'h00000086;
power_data[1591] = 32'h00000086;
power_data[1592] = 32'h00000086;
power_data[1593] = 32'h00000086;
power_data[1594] = 32'h00000086;
power_data[1595] = 32'h00000086;
power_data[1596] = 32'h00000086;
power_data[1597] = 32'h00000086;
power_data[1598] = 32'h00000086;
power_data[1599] = 32'h00000086;
power_data[1600] = 32'h00000086;
power_data[1601] = 32'h00000086;
power_data[1602] = 32'h00000086;
power_data[1603] = 32'h00000086;
power_data[1604] = 32'h00000086;
power_data[1605] = 32'h00000086;
power_data[1606] = 32'h00000086;
power_data[1607] = 32'h00000086;
power_data[1608] = 32'h00000086;
power_data[1609] = 32'h00000086;
power_data[1610] = 32'h00000086;
power_data[1611] = 32'h00000086;
power_data[1612] = 32'h00000086;
power_data[1613] = 32'h00000086;
power_data[1614] = 32'h00000086;
power_data[1615] = 32'h00000086;
power_data[1616] = 32'h00000086;
power_data[1617] = 32'h00000086;
power_data[1618] = 32'h00000086;
power_data[1619] = 32'h00000086;
power_data[1620] = 32'h00000086;
power_data[1621] = 32'h00000086;
power_data[1622] = 32'h00000086;
power_data[1623] = 32'h00000086;
power_data[1624] = 32'h00000086;
power_data[1625] = 32'h00000086;
power_data[1626] = 32'h00000086;
power_data[1627] = 32'h00000086;
power_data[1628] = 32'h00000086;
power_data[1629] = 32'h00000086;
power_data[1630] = 32'h00000086;
power_data[1631] = 32'h00000086;
power_data[1632] = 32'h00000086;
power_data[1633] = 32'h00000086;
power_data[1634] = 32'h00000086;
power_data[1635] = 32'h00000086;
power_data[1636] = 32'h00000086;
power_data[1637] = 32'h00000086;
power_data[1638] = 32'h00000086;
power_data[1639] = 32'h00000086;
power_data[1640] = 32'h00000086;
power_data[1641] = 32'h00000086;
power_data[1642] = 32'h00000086;
power_data[1643] = 32'h00000086;
power_data[1644] = 32'h00000086;
power_data[1645] = 32'h00000086;
power_data[1646] = 32'h00000086;
power_data[1647] = 32'h00000086;
power_data[1648] = 32'h00000086;
power_data[1649] = 32'h00000086;
power_data[1650] = 32'h00000086;
power_data[1651] = 32'h00000086;
power_data[1652] = 32'h00000086;
power_data[1653] = 32'h00000086;
power_data[1654] = 32'h00000086;
power_data[1655] = 32'h00000086;
power_data[1656] = 32'h00000086;
power_data[1657] = 32'h00000086;
power_data[1658] = 32'h00000086;
power_data[1659] = 32'h00000086;
power_data[1660] = 32'h00000086;
power_data[1661] = 32'h00000086;
power_data[1662] = 32'h00000086;
power_data[1663] = 32'h00000086;
power_data[1664] = 32'h00000086;
power_data[1665] = 32'h00000086;
power_data[1666] = 32'h00000086;
power_data[1667] = 32'h00000086;
power_data[1668] = 32'h00000086;
power_data[1669] = 32'h00000086;
power_data[1670] = 32'h00000086;
power_data[1671] = 32'h00000086;
power_data[1672] = 32'h00000086;
power_data[1673] = 32'h00000086;
power_data[1674] = 32'h00000086;
power_data[1675] = 32'h00000086;
power_data[1676] = 32'h00000086;
power_data[1677] = 32'h00000086;
power_data[1678] = 32'h00000086;
power_data[1679] = 32'h00000086;
power_data[1680] = 32'h00000086;
power_data[1681] = 32'h00000086;
power_data[1682] = 32'h00000086;
power_data[1683] = 32'h00000086;
power_data[1684] = 32'h00000086;
power_data[1685] = 32'h00000086;
power_data[1686] = 32'h00000086;
power_data[1687] = 32'h00000086;
power_data[1688] = 32'h00000086;
power_data[1689] = 32'h00000086;
power_data[1690] = 32'h00000086;
power_data[1691] = 32'h00000082;
power_data[1692] = 32'h00000069;
power_data[1693] = 32'h00000069;
power_data[1694] = 32'h00000069;
power_data[1695] = 32'h00000069;
power_data[1696] = 32'h00000069;
power_data[1697] = 32'h00000069;
power_data[1698] = 32'h00000069;
power_data[1699] = 32'h00000069;
power_data[1700] = 32'h00000069;
power_data[1701] = 32'h00000069;
power_data[1702] = 32'h00000069;
power_data[1703] = 32'h00000069;
power_data[1704] = 32'h00000069;
power_data[1705] = 32'h00000069;
power_data[1706] = 32'h00000069;
power_data[1707] = 32'h00000069;
power_data[1708] = 32'h00000069;
power_data[1709] = 32'h00000069;
power_data[1710] = 32'h00000069;
power_data[1711] = 32'h00000069;
power_data[1712] = 32'h00000069;
power_data[1713] = 32'h00000069;
power_data[1714] = 32'h00000069;
power_data[1715] = 32'h00000069;
power_data[1716] = 32'h00000069;
power_data[1717] = 32'h00000069;
power_data[1718] = 32'h00000069;
power_data[1719] = 32'h00000069;
power_data[1720] = 32'h00000069;
power_data[1721] = 32'h00000069;
power_data[1722] = 32'h00000069;
power_data[1723] = 32'h00000069;
power_data[1724] = 32'h00000069;
power_data[1725] = 32'h00000069;
power_data[1726] = 32'h00000069;
power_data[1727] = 32'h00000069;
power_data[1728] = 32'h00000069;
power_data[1729] = 32'h00000069;
power_data[1730] = 32'h00000069;
power_data[1731] = 32'h00000069;
power_data[1732] = 32'h00000069;
power_data[1733] = 32'h00000069;
power_data[1734] = 32'h00000069;
power_data[1735] = 32'h00000069;
power_data[1736] = 32'h00000069;
power_data[1737] = 32'h00000069;
power_data[1738] = 32'h00000069;
power_data[1739] = 32'h00000069;
power_data[1740] = 32'h00000069;
power_data[1741] = 32'h00000069;
power_data[1742] = 32'h00000069;
power_data[1743] = 32'h00000069;
power_data[1744] = 32'h00000069;
power_data[1745] = 32'h00000069;
power_data[1746] = 32'h00000069;
power_data[1747] = 32'h00000069;
power_data[1748] = 32'h00000069;
power_data[1749] = 32'h00000069;
power_data[1750] = 32'h00000069;
power_data[1751] = 32'h00000069;
power_data[1752] = 32'h00000069;
power_data[1753] = 32'h00000069;
power_data[1754] = 32'h00000069;
power_data[1755] = 32'h00000069;
power_data[1756] = 32'h00000069;
power_data[1757] = 32'h00000069;
power_data[1758] = 32'h00000069;
power_data[1759] = 32'h00000069;
power_data[1760] = 32'h00000069;
power_data[1761] = 32'h00000069;
power_data[1762] = 32'h0000077d;
power_data[1763] = 32'h00000942;
power_data[1764] = 32'h00000942;
power_data[1765] = 32'h00000942;
power_data[1766] = 32'h00000942;
power_data[1767] = 32'h00000942;
power_data[1768] = 32'h00000942;
power_data[1769] = 32'h00000942;
power_data[1770] = 32'h00000942;
power_data[1771] = 32'h00000942;
power_data[1772] = 32'h00000942;
power_data[1773] = 32'h00000942;
power_data[1774] = 32'h00000942;
power_data[1775] = 32'h00000942;
power_data[1776] = 32'h00000942;
power_data[1777] = 32'h00000942;
power_data[1778] = 32'h00000942;
power_data[1779] = 32'h00000942;
power_data[1780] = 32'h00000942;
power_data[1781] = 32'h00000942;
power_data[1782] = 32'h00000942;
power_data[1783] = 32'h00000942;
power_data[1784] = 32'h00000942;
power_data[1785] = 32'h00000942;
power_data[1786] = 32'h00000942;
power_data[1787] = 32'h00000942;
power_data[1788] = 32'h00000942;
power_data[1789] = 32'h00000942;
power_data[1790] = 32'h00000942;
power_data[1791] = 32'h00000232;
power_data[1792] = 32'h00000232;
power_data[1793] = 32'h00000232;
power_data[1794] = 32'h00000232;
power_data[1795] = 32'h00000232;
power_data[1796] = 32'h00000232;
power_data[1797] = 32'h00000232;
power_data[1798] = 32'h00000232;
power_data[1799] = 32'h00000232;
power_data[1800] = 32'h00000232;
power_data[1801] = 32'h00000232;
power_data[1802] = 32'h00000232;
power_data[1803] = 32'h00000232;
power_data[1804] = 32'h00000232;
power_data[1805] = 32'h00000232;
power_data[1806] = 32'h00000232;
power_data[1807] = 32'h00000232;
power_data[1808] = 32'h00000232;
power_data[1809] = 32'h00000232;
power_data[1810] = 32'h00000232;
power_data[1811] = 32'h00000232;
power_data[1812] = 32'h00000232;
power_data[1813] = 32'h00000232;
power_data[1814] = 32'h00000232;
power_data[1815] = 32'h00000232;
power_data[1816] = 32'h00000232;
power_data[1817] = 32'h00000232;
power_data[1818] = 32'h00000232;
power_data[1819] = 32'h00000232;
power_data[1820] = 32'h00000232;
power_data[1821] = 32'h00000232;
power_data[1822] = 32'h00000232;
power_data[1823] = 32'h00000232;
power_data[1824] = 32'h00000232;
power_data[1825] = 32'h00000232;
power_data[1826] = 32'h00000232;
power_data[1827] = 32'h00000232;
power_data[1828] = 32'h00000232;
power_data[1829] = 32'h00000232;
power_data[1830] = 32'h00000232;
power_data[1831] = 32'h00000232;
power_data[1832] = 32'h000013d3;
power_data[1833] = 32'h00002e41;
power_data[1834] = 32'h00002e41;
power_data[1835] = 32'h00002e41;
power_data[1836] = 32'h00002e41;
power_data[1837] = 32'h00002e41;
power_data[1838] = 32'h00002e41;
power_data[1839] = 32'h00002e41;
power_data[1840] = 32'h00002e41;
power_data[1841] = 32'h00002e41;
power_data[1842] = 32'h00002e41;
power_data[1843] = 32'h00002e41;
power_data[1844] = 32'h00002e41;
power_data[1845] = 32'h00002e41;
power_data[1846] = 32'h00002e41;
power_data[1847] = 32'h00002e41;
power_data[1848] = 32'h00002e41;
power_data[1849] = 32'h00002e41;
power_data[1850] = 32'h00002e41;
power_data[1851] = 32'h00002e41;
power_data[1852] = 32'h00002e41;
power_data[1853] = 32'h00002e41;
power_data[1854] = 32'h00002e41;
power_data[1855] = 32'h00002e41;
power_data[1856] = 32'h00002e41;
power_data[1857] = 32'h00002e41;
power_data[1858] = 32'h00002e41;
power_data[1859] = 32'h00002e41;
power_data[1860] = 32'h00002e41;
power_data[1861] = 32'h00002e41;
power_data[1862] = 32'h00002e41;
power_data[1863] = 32'h00002e41;
power_data[1864] = 32'h00002e41;
power_data[1865] = 32'h00002e41;
power_data[1866] = 32'h00002e41;
power_data[1867] = 32'h00002e41;
power_data[1868] = 32'h00002e41;
power_data[1869] = 32'h00002e41;
power_data[1870] = 32'h00002e41;
power_data[1871] = 32'h00002e41;
power_data[1872] = 32'h00002e41;
power_data[1873] = 32'h00002e41;
power_data[1874] = 32'h00002e41;
power_data[1875] = 32'h00002e41;
power_data[1876] = 32'h00002e41;
power_data[1877] = 32'h00002e41;
power_data[1878] = 32'h00002e41;
power_data[1879] = 32'h00002e41;
power_data[1880] = 32'h00002e41;
power_data[1881] = 32'h00002e41;
power_data[1882] = 32'h00002e41;
power_data[1883] = 32'h00002e41;
power_data[1884] = 32'h00002e41;
power_data[1885] = 32'h00002e41;
power_data[1886] = 32'h00002e41;
power_data[1887] = 32'h00002e41;
power_data[1888] = 32'h00002e41;
power_data[1889] = 32'h00002e41;
power_data[1890] = 32'h000009ab;
power_data[1891] = 32'h00000086;
power_data[1892] = 32'h00000086;
power_data[1893] = 32'h00000086;
power_data[1894] = 32'h00000086;
power_data[1895] = 32'h00000086;
power_data[1896] = 32'h00000086;
power_data[1897] = 32'h00000086;
power_data[1898] = 32'h00000086;
power_data[1899] = 32'h00000086;
power_data[1900] = 32'h00000086;
power_data[1901] = 32'h00000086;
power_data[1902] = 32'h00000086;
power_data[1903] = 32'h00000086;
power_data[1904] = 32'h00000086;
power_data[1905] = 32'h00000086;
power_data[1906] = 32'h00000086;
power_data[1907] = 32'h00000086;
power_data[1908] = 32'h00000086;
power_data[1909] = 32'h00000086;
power_data[1910] = 32'h00000086;
power_data[1911] = 32'h00000086;
power_data[1912] = 32'h00000086;
power_data[1913] = 32'h00000086;
power_data[1914] = 32'h00000086;
power_data[1915] = 32'h00000086;
power_data[1916] = 32'h00000086;
power_data[1917] = 32'h00000086;
power_data[1918] = 32'h00000086;
power_data[1919] = 32'h00000086;
power_data[1920] = 32'h00000086;
power_data[1921] = 32'h00000086;
power_data[1922] = 32'h00000086;
power_data[1923] = 32'h00000086;
power_data[1924] = 32'h00000086;
power_data[1925] = 32'h00000086;
power_data[1926] = 32'h00000086;
power_data[1927] = 32'h00000086;
power_data[1928] = 32'h00000086;
power_data[1929] = 32'h00000086;
power_data[1930] = 32'h00000086;
power_data[1931] = 32'h00000086;
power_data[1932] = 32'h00000086;
power_data[1933] = 32'h00000086;
power_data[1934] = 32'h00000086;
power_data[1935] = 32'h00000086;
power_data[1936] = 32'h00000086;
power_data[1937] = 32'h00000086;
power_data[1938] = 32'h00000086;
power_data[1939] = 32'h00000086;
power_data[1940] = 32'h00000086;
power_data[1941] = 32'h00000086;
power_data[1942] = 32'h00000086;
power_data[1943] = 32'h00000086;
power_data[1944] = 32'h00000086;
power_data[1945] = 32'h00000086;
power_data[1946] = 32'h00000086;
power_data[1947] = 32'h00000086;
power_data[1948] = 32'h00000086;
power_data[1949] = 32'h00000086;
power_data[1950] = 32'h00000086;
power_data[1951] = 32'h00000086;
power_data[1952] = 32'h00000086;
power_data[1953] = 32'h00000086;
power_data[1954] = 32'h00000086;
power_data[1955] = 32'h00000086;
power_data[1956] = 32'h00000086;
power_data[1957] = 32'h00000086;
power_data[1958] = 32'h00000086;
power_data[1959] = 32'h00000086;
power_data[1960] = 32'h00000086;
power_data[1961] = 32'h00000086;
power_data[1962] = 32'h00000086;
power_data[1963] = 32'h00000086;
power_data[1964] = 32'h00000086;
power_data[1965] = 32'h00000086;
power_data[1966] = 32'h00000086;
power_data[1967] = 32'h00000086;
power_data[1968] = 32'h00000086;
power_data[1969] = 32'h00000086;
power_data[1970] = 32'h00000086;
power_data[1971] = 32'h00000086;
power_data[1972] = 32'h00000086;
power_data[1973] = 32'h00000086;
power_data[1974] = 32'h00000086;
power_data[1975] = 32'h00000086;
power_data[1976] = 32'h00000086;
power_data[1977] = 32'h00000086;
power_data[1978] = 32'h00000086;
power_data[1979] = 32'h00000086;
power_data[1980] = 32'h00000086;
power_data[1981] = 32'h00000086;
power_data[1982] = 32'h00000086;
power_data[1983] = 32'h00000086;
power_data[1984] = 32'h00000086;
power_data[1985] = 32'h00000086;
power_data[1986] = 32'h00000086;
power_data[1987] = 32'h00000086;
power_data[1988] = 32'h00000086;
power_data[1989] = 32'h00000086;
power_data[1990] = 32'h00000086;
power_data[1991] = 32'h00000086;
power_data[1992] = 32'h00000086;
power_data[1993] = 32'h00000086;
power_data[1994] = 32'h00000086;
power_data[1995] = 32'h00000086;
power_data[1996] = 32'h00000086;
power_data[1997] = 32'h00000086;
power_data[1998] = 32'h00000086;
power_data[1999] = 32'h00000086;
power_data[2000] = 32'h00000086;
power_data[2001] = 32'h00000086;
power_data[2002] = 32'h00000086;
power_data[2003] = 32'h00000086;
power_data[2004] = 32'h00000086;
power_data[2005] = 32'h00000086;
power_data[2006] = 32'h00000086;
power_data[2007] = 32'h00000086;
power_data[2008] = 32'h00000086;
power_data[2009] = 32'h00000086;
power_data[2010] = 32'h00000086;
power_data[2011] = 32'h00000086;
power_data[2012] = 32'h00000086;
power_data[2013] = 32'h00000086;
power_data[2014] = 32'h00000086;
power_data[2015] = 32'h00000086;
power_data[2016] = 32'h00000086;
power_data[2017] = 32'h00000086;
power_data[2018] = 32'h00000086;
power_data[2019] = 32'h00000086;
power_data[2020] = 32'h00000086;
power_data[2021] = 32'h00000086;
power_data[2022] = 32'h00000086;
power_data[2023] = 32'h00000086;
power_data[2024] = 32'h00000086;
power_data[2025] = 32'h00000086;
power_data[2026] = 32'h00000086;
power_data[2027] = 32'h00000086;
power_data[2028] = 32'h00000086;
power_data[2029] = 32'h00000086;
power_data[2030] = 32'h00000086;
power_data[2031] = 32'h00000086;
power_data[2032] = 32'h00000086;
power_data[2033] = 32'h00000086;
power_data[2034] = 32'h00000086;
power_data[2035] = 32'h00000086;
power_data[2036] = 32'h00000086;
power_data[2037] = 32'h00000086;
power_data[2038] = 32'h00000086;
power_data[2039] = 32'h00000086;
power_data[2040] = 32'h00000086;
power_data[2041] = 32'h00000086;
power_data[2042] = 32'h00000086;
power_data[2043] = 32'h00000086;
power_data[2044] = 32'h00000086;
power_data[2045] = 32'h00000086;
power_data[2046] = 32'h00000086;
power_data[2047] = 32'h00000086;
power_data[2048] = 32'h00000086;
power_data[2049] = 32'h00000086;
power_data[2050] = 32'h00000086;
power_data[2051] = 32'h00000086;
power_data[2052] = 32'h00000086;
power_data[2053] = 32'h00000086;
power_data[2054] = 32'h00000086;
power_data[2055] = 32'h00000086;
power_data[2056] = 32'h00000086;
power_data[2057] = 32'h00000086;
power_data[2058] = 32'h00000086;
power_data[2059] = 32'h00000086;
power_data[2060] = 32'h00000086;
power_data[2061] = 32'h00000086;
power_data[2062] = 32'h00000086;
power_data[2063] = 32'h00000086;
power_data[2064] = 32'h00000086;
power_data[2065] = 32'h00000086;
power_data[2066] = 32'h00000086;
power_data[2067] = 32'h00000086;
power_data[2068] = 32'h00000086;
power_data[2069] = 32'h00000086;
power_data[2070] = 32'h00000086;
power_data[2071] = 32'h00000086;
power_data[2072] = 32'h00000086;
power_data[2073] = 32'h00000086;
power_data[2074] = 32'h00000086;
power_data[2075] = 32'h00000086;
power_data[2076] = 32'h00000086;
power_data[2077] = 32'h00000086;
power_data[2078] = 32'h00000086;
power_data[2079] = 32'h00000086;
power_data[2080] = 32'h00000086;
power_data[2081] = 32'h00000086;
power_data[2082] = 32'h00000086;
power_data[2083] = 32'h00000086;
power_data[2084] = 32'h00000086;
power_data[2085] = 32'h00000086;
power_data[2086] = 32'h00000086;
power_data[2087] = 32'h00000086;
power_data[2088] = 32'h00000086;
power_data[2089] = 32'h00000086;
power_data[2090] = 32'h00000086;
power_data[2091] = 32'h00000086;
power_data[2092] = 32'h00000086;
power_data[2093] = 32'h00000086;
power_data[2094] = 32'h00000086;
power_data[2095] = 32'h00000086;
power_data[2096] = 32'h00000086;
power_data[2097] = 32'h00000086;
power_data[2098] = 32'h00000086;
power_data[2099] = 32'h00000086;
power_data[2100] = 32'h00000086;
power_data[2101] = 32'h00000086;
power_data[2102] = 32'h00000086;
power_data[2103] = 32'h00000086;
power_data[2104] = 32'h00000086;
power_data[2105] = 32'h00000086;
power_data[2106] = 32'h00000086;
power_data[2107] = 32'h00000086;
power_data[2108] = 32'h00000086;
power_data[2109] = 32'h00000086;
power_data[2110] = 32'h00000086;
power_data[2111] = 32'h00000086;
power_data[2112] = 32'h00000086;
power_data[2113] = 32'h00000086;
power_data[2114] = 32'h00000086;
power_data[2115] = 32'h00000086;
power_data[2116] = 32'h00000086;
power_data[2117] = 32'h00000086;
power_data[2118] = 32'h00000086;
power_data[2119] = 32'h00000086;
power_data[2120] = 32'h00000086;
power_data[2121] = 32'h00000086;
power_data[2122] = 32'h00000086;
power_data[2123] = 32'h00000086;
power_data[2124] = 32'h00000086;
power_data[2125] = 32'h00000086;
power_data[2126] = 32'h00000086;
power_data[2127] = 32'h00000086;
power_data[2128] = 32'h00000086;
power_data[2129] = 32'h00000086;
power_data[2130] = 32'h00000086;
power_data[2131] = 32'h00000086;
power_data[2132] = 32'h00000086;
power_data[2133] = 32'h00000086;
power_data[2134] = 32'h00000086;
power_data[2135] = 32'h00000086;
power_data[2136] = 32'h00000086;
power_data[2137] = 32'h00000086;
power_data[2138] = 32'h00000086;
power_data[2139] = 32'h00000086;
power_data[2140] = 32'h00000086;
power_data[2141] = 32'h00000086;
power_data[2142] = 32'h00000086;
power_data[2143] = 32'h00000086;
power_data[2144] = 32'h00000086;
power_data[2145] = 32'h00000086;
power_data[2146] = 32'h00000086;
power_data[2147] = 32'h00000086;
power_data[2148] = 32'h00000086;
power_data[2149] = 32'h00000086;
power_data[2150] = 32'h00000086;
power_data[2151] = 32'h00000086;
power_data[2152] = 32'h00000086;
power_data[2153] = 32'h00000086;
power_data[2154] = 32'h00000086;
power_data[2155] = 32'h00000086;
power_data[2156] = 32'h00000086;
power_data[2157] = 32'h00000086;
power_data[2158] = 32'h00000086;
power_data[2159] = 32'h00000086;
power_data[2160] = 32'h00000086;
power_data[2161] = 32'h00000086;
power_data[2162] = 32'h00000086;
power_data[2163] = 32'h00000086;
power_data[2164] = 32'h00000086;
power_data[2165] = 32'h00000086;
power_data[2166] = 32'h00000086;
power_data[2167] = 32'h00000086;
power_data[2168] = 32'h00000086;
power_data[2169] = 32'h00000086;
power_data[2170] = 32'h00000086;
power_data[2171] = 32'h00000086;
power_data[2172] = 32'h00000086;
power_data[2173] = 32'h00000086;
power_data[2174] = 32'h00000086;
power_data[2175] = 32'h00000086;
power_data[2176] = 32'h00000086;
power_data[2177] = 32'h00000086;
power_data[2178] = 32'h00000086;
power_data[2179] = 32'h00000086;
power_data[2180] = 32'h00000086;
power_data[2181] = 32'h00000086;
power_data[2182] = 32'h00000086;
power_data[2183] = 32'h00000086;
power_data[2184] = 32'h00000086;
power_data[2185] = 32'h00000086;
power_data[2186] = 32'h00000086;
power_data[2187] = 32'h00000086;
power_data[2188] = 32'h00000086;
power_data[2189] = 32'h00000086;
power_data[2190] = 32'h00000086;
power_data[2191] = 32'h00000086;
power_data[2192] = 32'h00000086;
power_data[2193] = 32'h00000086;
power_data[2194] = 32'h00000086;
power_data[2195] = 32'h00000086;
power_data[2196] = 32'h00000086;
power_data[2197] = 32'h00000086;
power_data[2198] = 32'h00000086;
power_data[2199] = 32'h00000086;
power_data[2200] = 32'h00000086;
power_data[2201] = 32'h00000086;
power_data[2202] = 32'h00000086;
power_data[2203] = 32'h00000082;
power_data[2204] = 32'h00000069;
power_data[2205] = 32'h00000069;
power_data[2206] = 32'h00000069;
power_data[2207] = 32'h00000069;
power_data[2208] = 32'h00000069;
power_data[2209] = 32'h00000069;
power_data[2210] = 32'h00000069;
power_data[2211] = 32'h00000069;
power_data[2212] = 32'h00000069;
power_data[2213] = 32'h00000069;
power_data[2214] = 32'h00000069;
power_data[2215] = 32'h00000069;
power_data[2216] = 32'h00000069;
power_data[2217] = 32'h00000069;
power_data[2218] = 32'h00000069;
power_data[2219] = 32'h00000069;
power_data[2220] = 32'h00000069;
power_data[2221] = 32'h00000069;
power_data[2222] = 32'h00000069;
power_data[2223] = 32'h00000069;
power_data[2224] = 32'h00000069;
power_data[2225] = 32'h00000069;
power_data[2226] = 32'h00000069;
power_data[2227] = 32'h00000069;
power_data[2228] = 32'h00000069;
power_data[2229] = 32'h00000069;
power_data[2230] = 32'h00000069;
power_data[2231] = 32'h00000069;
power_data[2232] = 32'h00000069;
power_data[2233] = 32'h00000069;
power_data[2234] = 32'h00000069;
power_data[2235] = 32'h00000069;
power_data[2236] = 32'h00000069;
power_data[2237] = 32'h00000069;
power_data[2238] = 32'h00000069;
power_data[2239] = 32'h00000069;
power_data[2240] = 32'h00000069;
power_data[2241] = 32'h00000069;
power_data[2242] = 32'h00000069;
power_data[2243] = 32'h00000069;
power_data[2244] = 32'h00000069;
power_data[2245] = 32'h00000069;
power_data[2246] = 32'h00000069;
power_data[2247] = 32'h00000069;
power_data[2248] = 32'h00000069;
power_data[2249] = 32'h00000069;
power_data[2250] = 32'h00000069;
power_data[2251] = 32'h00000069;
power_data[2252] = 32'h00000069;
power_data[2253] = 32'h00000069;
power_data[2254] = 32'h00000069;
power_data[2255] = 32'h00000069;
power_data[2256] = 32'h00000069;
power_data[2257] = 32'h00000069;
power_data[2258] = 32'h00000069;
power_data[2259] = 32'h00000069;
power_data[2260] = 32'h00000069;
power_data[2261] = 32'h00000069;
power_data[2262] = 32'h00000069;
power_data[2263] = 32'h00000069;
power_data[2264] = 32'h00000069;
power_data[2265] = 32'h00000069;
power_data[2266] = 32'h00000069;
power_data[2267] = 32'h00000069;
power_data[2268] = 32'h00000069;
power_data[2269] = 32'h00000069;
power_data[2270] = 32'h00000069;
power_data[2271] = 32'h00000069;
power_data[2272] = 32'h00000069;
power_data[2273] = 32'h00000069;
power_data[2274] = 32'h0000077d;
power_data[2275] = 32'h00000942;
power_data[2276] = 32'h00000942;
power_data[2277] = 32'h00000942;
power_data[2278] = 32'h00000942;
power_data[2279] = 32'h00000942;
power_data[2280] = 32'h00000942;
power_data[2281] = 32'h00000942;
power_data[2282] = 32'h00000942;
power_data[2283] = 32'h00000942;
power_data[2284] = 32'h00000942;
power_data[2285] = 32'h00000942;
power_data[2286] = 32'h00000942;
power_data[2287] = 32'h00000942;
power_data[2288] = 32'h00000942;
power_data[2289] = 32'h00000942;
power_data[2290] = 32'h00000942;
power_data[2291] = 32'h00000942;
power_data[2292] = 32'h00000942;
power_data[2293] = 32'h00000942;
power_data[2294] = 32'h00000942;
power_data[2295] = 32'h00000942;
power_data[2296] = 32'h00000942;
power_data[2297] = 32'h00000942;
power_data[2298] = 32'h00000942;
power_data[2299] = 32'h00000942;
power_data[2300] = 32'h00000942;
power_data[2301] = 32'h00000942;
power_data[2302] = 32'h00000942;
power_data[2303] = 32'h00000232;
power_data[2304] = 32'h00000232;
power_data[2305] = 32'h00000232;
power_data[2306] = 32'h00000232;
power_data[2307] = 32'h00000232;
power_data[2308] = 32'h00000232;
power_data[2309] = 32'h00000232;
power_data[2310] = 32'h00000232;
power_data[2311] = 32'h00000232;
power_data[2312] = 32'h00000232;
power_data[2313] = 32'h00000232;
power_data[2314] = 32'h00000232;
power_data[2315] = 32'h00000232;
power_data[2316] = 32'h00000232;
power_data[2317] = 32'h00000232;
power_data[2318] = 32'h00000232;
power_data[2319] = 32'h00000232;
power_data[2320] = 32'h00000232;
power_data[2321] = 32'h00000232;
power_data[2322] = 32'h00000232;
power_data[2323] = 32'h00000232;
power_data[2324] = 32'h00000232;
power_data[2325] = 32'h00000232;
power_data[2326] = 32'h00000232;
power_data[2327] = 32'h00000232;
power_data[2328] = 32'h00000232;
power_data[2329] = 32'h00000232;
power_data[2330] = 32'h00000232;
power_data[2331] = 32'h00000232;
power_data[2332] = 32'h00000232;
power_data[2333] = 32'h00000232;
power_data[2334] = 32'h00000232;
power_data[2335] = 32'h00000232;
power_data[2336] = 32'h00000232;
power_data[2337] = 32'h00000232;
power_data[2338] = 32'h00000232;
power_data[2339] = 32'h00000232;
power_data[2340] = 32'h00000232;
power_data[2341] = 32'h00000232;
power_data[2342] = 32'h00000232;
power_data[2343] = 32'h00000232;
power_data[2344] = 32'h000013d3;
power_data[2345] = 32'h00002e41;
power_data[2346] = 32'h00002e41;
power_data[2347] = 32'h00002e41;
power_data[2348] = 32'h00002e41;
power_data[2349] = 32'h00002e41;
power_data[2350] = 32'h00002e41;
power_data[2351] = 32'h00002e41;
power_data[2352] = 32'h00002e41;
power_data[2353] = 32'h00002e41;
power_data[2354] = 32'h00002e41;
power_data[2355] = 32'h00002e41;
power_data[2356] = 32'h00002e41;
power_data[2357] = 32'h00002e41;
power_data[2358] = 32'h00002e41;
power_data[2359] = 32'h00002e41;
power_data[2360] = 32'h00002e41;
power_data[2361] = 32'h00002e41;
power_data[2362] = 32'h00002e41;
power_data[2363] = 32'h00002e41;
power_data[2364] = 32'h00002e41;
power_data[2365] = 32'h00002e41;
power_data[2366] = 32'h00002e41;
power_data[2367] = 32'h00002e41;
power_data[2368] = 32'h00002e41;
power_data[2369] = 32'h00002e41;
power_data[2370] = 32'h00002e41;
power_data[2371] = 32'h00002e41;
power_data[2372] = 32'h00002e41;
power_data[2373] = 32'h00002e41;
power_data[2374] = 32'h00002e41;
power_data[2375] = 32'h00002e41;
power_data[2376] = 32'h00002e41;
power_data[2377] = 32'h00002e41;
power_data[2378] = 32'h00002e41;
power_data[2379] = 32'h00002e41;
power_data[2380] = 32'h00002e41;
power_data[2381] = 32'h00002e41;
power_data[2382] = 32'h00002e41;
power_data[2383] = 32'h00002e41;
power_data[2384] = 32'h00002e41;
power_data[2385] = 32'h00002e41;
power_data[2386] = 32'h00002e41;
power_data[2387] = 32'h00002e41;
power_data[2388] = 32'h00002e41;
power_data[2389] = 32'h00002e41;
power_data[2390] = 32'h00002e41;
power_data[2391] = 32'h00002e41;
power_data[2392] = 32'h00002e41;
power_data[2393] = 32'h00002e41;
power_data[2394] = 32'h00002e41;
power_data[2395] = 32'h00002e41;
power_data[2396] = 32'h00002e41;
power_data[2397] = 32'h00002e41;
power_data[2398] = 32'h00002e41;
power_data[2399] = 32'h00002e41;
power_data[2400] = 32'h00002e41;
power_data[2401] = 32'h00002e41;
power_data[2402] = 32'h000009ab;
power_data[2403] = 32'h00000086;
power_data[2404] = 32'h00000086;
power_data[2405] = 32'h00000086;
power_data[2406] = 32'h00000086;
power_data[2407] = 32'h00000086;
power_data[2408] = 32'h00000086;
power_data[2409] = 32'h00000086;
power_data[2410] = 32'h00000086;
power_data[2411] = 32'h00000086;
power_data[2412] = 32'h00000086;
power_data[2413] = 32'h00000086;
power_data[2414] = 32'h00000086;
power_data[2415] = 32'h00000086;
power_data[2416] = 32'h00000086;
power_data[2417] = 32'h00000086;
power_data[2418] = 32'h00000086;
power_data[2419] = 32'h00000086;
power_data[2420] = 32'h00000086;
power_data[2421] = 32'h00000086;
power_data[2422] = 32'h00000086;
power_data[2423] = 32'h00000086;
power_data[2424] = 32'h00000086;
power_data[2425] = 32'h00000086;
power_data[2426] = 32'h00000086;
power_data[2427] = 32'h00000086;
power_data[2428] = 32'h00000086;
power_data[2429] = 32'h00000086;
power_data[2430] = 32'h00000086;
power_data[2431] = 32'h00000086;
power_data[2432] = 32'h00000086;
power_data[2433] = 32'h00000086;
power_data[2434] = 32'h00000086;
power_data[2435] = 32'h00000086;
power_data[2436] = 32'h00000086;
power_data[2437] = 32'h00000086;
power_data[2438] = 32'h00000086;
power_data[2439] = 32'h00000086;
power_data[2440] = 32'h00000086;
power_data[2441] = 32'h00000086;
power_data[2442] = 32'h00000086;
power_data[2443] = 32'h00000086;
power_data[2444] = 32'h00000086;
power_data[2445] = 32'h00000086;
power_data[2446] = 32'h00000086;
power_data[2447] = 32'h00000086;
power_data[2448] = 32'h00000086;
power_data[2449] = 32'h00000086;
power_data[2450] = 32'h00000086;
power_data[2451] = 32'h00000086;
power_data[2452] = 32'h00000086;
power_data[2453] = 32'h00000086;
power_data[2454] = 32'h00000086;
power_data[2455] = 32'h00000086;
power_data[2456] = 32'h00000086;
power_data[2457] = 32'h00000086;
power_data[2458] = 32'h00000086;
power_data[2459] = 32'h00000086;
power_data[2460] = 32'h00000086;
power_data[2461] = 32'h00000086;
power_data[2462] = 32'h00000086;
power_data[2463] = 32'h00000086;
power_data[2464] = 32'h00000086;
power_data[2465] = 32'h00000086;
power_data[2466] = 32'h00000086;
power_data[2467] = 32'h00000086;
power_data[2468] = 32'h00000086;
power_data[2469] = 32'h00000086;
power_data[2470] = 32'h00000086;
power_data[2471] = 32'h00000086;
power_data[2472] = 32'h00000086;
power_data[2473] = 32'h00000086;
power_data[2474] = 32'h00000086;
power_data[2475] = 32'h00000086;
power_data[2476] = 32'h00000086;
power_data[2477] = 32'h00000086;
power_data[2478] = 32'h00000086;
power_data[2479] = 32'h00000086;
power_data[2480] = 32'h00000086;
power_data[2481] = 32'h00000086;
power_data[2482] = 32'h00000086;
power_data[2483] = 32'h00000086;
power_data[2484] = 32'h00000086;
power_data[2485] = 32'h00000086;
power_data[2486] = 32'h00000086;
power_data[2487] = 32'h00000086;
power_data[2488] = 32'h00000086;
power_data[2489] = 32'h00000086;
power_data[2490] = 32'h00000086;
power_data[2491] = 32'h00000086;
power_data[2492] = 32'h00000086;
power_data[2493] = 32'h00000086;
power_data[2494] = 32'h00000086;
power_data[2495] = 32'h00000086;
power_data[2496] = 32'h00000086;
power_data[2497] = 32'h00000086;
power_data[2498] = 32'h00000086;
power_data[2499] = 32'h00000086;
power_data[2500] = 32'h00000086;
power_data[2501] = 32'h00000086;
power_data[2502] = 32'h00000086;
power_data[2503] = 32'h00000086;
power_data[2504] = 32'h00000086;
power_data[2505] = 32'h00000086;
power_data[2506] = 32'h00000086;
power_data[2507] = 32'h00000086;
power_data[2508] = 32'h00000086;
power_data[2509] = 32'h00000086;
power_data[2510] = 32'h00000086;
power_data[2511] = 32'h00000086;
power_data[2512] = 32'h00000086;
power_data[2513] = 32'h00000086;
power_data[2514] = 32'h00000086;
power_data[2515] = 32'h00000086;
power_data[2516] = 32'h00000086;
power_data[2517] = 32'h00000086;
power_data[2518] = 32'h00000086;
power_data[2519] = 32'h00000086;
power_data[2520] = 32'h00000086;
power_data[2521] = 32'h00000086;
power_data[2522] = 32'h00000086;
power_data[2523] = 32'h00000086;
power_data[2524] = 32'h00000086;
power_data[2525] = 32'h00000086;
power_data[2526] = 32'h00000086;
power_data[2527] = 32'h00000086;
power_data[2528] = 32'h00000086;
power_data[2529] = 32'h00000086;
power_data[2530] = 32'h00000086;
power_data[2531] = 32'h00000086;
power_data[2532] = 32'h00000086;
power_data[2533] = 32'h00000086;
power_data[2534] = 32'h00000086;
power_data[2535] = 32'h00000086;
power_data[2536] = 32'h00000086;
power_data[2537] = 32'h00000086;
power_data[2538] = 32'h00000086;
power_data[2539] = 32'h00000086;
power_data[2540] = 32'h00000086;
power_data[2541] = 32'h00000086;
power_data[2542] = 32'h00000086;
power_data[2543] = 32'h00000086;
power_data[2544] = 32'h00000086;
power_data[2545] = 32'h00000086;
power_data[2546] = 32'h00000086;
power_data[2547] = 32'h00000086;
power_data[2548] = 32'h00000086;
power_data[2549] = 32'h00000086;
power_data[2550] = 32'h00000086;
power_data[2551] = 32'h00000086;
power_data[2552] = 32'h00000086;
power_data[2553] = 32'h00000086;
power_data[2554] = 32'h00000086;
power_data[2555] = 32'h00000086;
power_data[2556] = 32'h00000086;
power_data[2557] = 32'h00000086;
power_data[2558] = 32'h00000086;
power_data[2559] = 32'h00000086;
power_data[2560] = 32'h00000086;
power_data[2561] = 32'h00000086;
power_data[2562] = 32'h00000086;
power_data[2563] = 32'h00000086;
power_data[2564] = 32'h00000086;
power_data[2565] = 32'h00000086;
power_data[2566] = 32'h00000086;
power_data[2567] = 32'h00000086;
power_data[2568] = 32'h00000086;
power_data[2569] = 32'h00000086;
power_data[2570] = 32'h00000086;
power_data[2571] = 32'h00000086;
power_data[2572] = 32'h00000086;
power_data[2573] = 32'h00000086;
power_data[2574] = 32'h00000086;
power_data[2575] = 32'h00000086;
power_data[2576] = 32'h00000086;
power_data[2577] = 32'h00000086;
power_data[2578] = 32'h00000086;
power_data[2579] = 32'h00000086;
power_data[2580] = 32'h00000086;
power_data[2581] = 32'h00000086;
power_data[2582] = 32'h00000086;
power_data[2583] = 32'h00000086;
power_data[2584] = 32'h00000086;
power_data[2585] = 32'h00000086;
power_data[2586] = 32'h00000086;
power_data[2587] = 32'h00000086;
power_data[2588] = 32'h00000086;
power_data[2589] = 32'h00000086;
power_data[2590] = 32'h00000086;
power_data[2591] = 32'h00000086;
power_data[2592] = 32'h00000086;
power_data[2593] = 32'h00000086;
power_data[2594] = 32'h00000086;
power_data[2595] = 32'h00000086;
power_data[2596] = 32'h00000086;
power_data[2597] = 32'h00000086;
power_data[2598] = 32'h00000086;
power_data[2599] = 32'h00000086;
power_data[2600] = 32'h00000086;
power_data[2601] = 32'h00000086;
power_data[2602] = 32'h00000086;
power_data[2603] = 32'h00000086;
power_data[2604] = 32'h00000086;
power_data[2605] = 32'h00000086;
power_data[2606] = 32'h00000086;
power_data[2607] = 32'h00000086;
power_data[2608] = 32'h00000086;
power_data[2609] = 32'h00000086;
power_data[2610] = 32'h00000086;
power_data[2611] = 32'h00000086;
power_data[2612] = 32'h00000086;
power_data[2613] = 32'h00000086;
power_data[2614] = 32'h00000086;
power_data[2615] = 32'h00000086;
power_data[2616] = 32'h00000086;
power_data[2617] = 32'h00000086;
power_data[2618] = 32'h00000086;
power_data[2619] = 32'h00000086;
power_data[2620] = 32'h00000086;
power_data[2621] = 32'h00000086;
power_data[2622] = 32'h00000086;
power_data[2623] = 32'h00000086;
power_data[2624] = 32'h00000086;
power_data[2625] = 32'h00000086;
power_data[2626] = 32'h00000086;
power_data[2627] = 32'h00000086;
power_data[2628] = 32'h00000086;
power_data[2629] = 32'h00000086;
power_data[2630] = 32'h00000086;
power_data[2631] = 32'h00000086;
power_data[2632] = 32'h00000086;
power_data[2633] = 32'h00000086;
power_data[2634] = 32'h00000086;
power_data[2635] = 32'h00000086;
power_data[2636] = 32'h00000086;
power_data[2637] = 32'h00000086;
power_data[2638] = 32'h00000086;
power_data[2639] = 32'h00000086;
power_data[2640] = 32'h00000086;
power_data[2641] = 32'h00000086;
power_data[2642] = 32'h00000086;
power_data[2643] = 32'h00000086;
power_data[2644] = 32'h00000086;
power_data[2645] = 32'h00000086;
power_data[2646] = 32'h00000086;
power_data[2647] = 32'h00000086;
power_data[2648] = 32'h00000086;
power_data[2649] = 32'h00000086;
power_data[2650] = 32'h00000086;
power_data[2651] = 32'h00000086;
power_data[2652] = 32'h00000086;
power_data[2653] = 32'h00000086;
power_data[2654] = 32'h00000086;
power_data[2655] = 32'h00000086;
power_data[2656] = 32'h00000086;
power_data[2657] = 32'h00000086;
power_data[2658] = 32'h00000086;
power_data[2659] = 32'h00000086;
power_data[2660] = 32'h00000086;
power_data[2661] = 32'h00000086;
power_data[2662] = 32'h00000086;
power_data[2663] = 32'h00000086;
power_data[2664] = 32'h00000086;
power_data[2665] = 32'h00000086;
power_data[2666] = 32'h00000086;
power_data[2667] = 32'h00000086;
power_data[2668] = 32'h00000086;
power_data[2669] = 32'h00000086;
power_data[2670] = 32'h00000086;
power_data[2671] = 32'h00000086;
power_data[2672] = 32'h00000086;
power_data[2673] = 32'h00000086;
power_data[2674] = 32'h00000086;
power_data[2675] = 32'h00000086;
power_data[2676] = 32'h00000086;
power_data[2677] = 32'h00000086;
power_data[2678] = 32'h00000086;
power_data[2679] = 32'h00000086;
power_data[2680] = 32'h00000086;
power_data[2681] = 32'h00000086;
power_data[2682] = 32'h00000086;
power_data[2683] = 32'h00000086;
power_data[2684] = 32'h00000086;
power_data[2685] = 32'h00000086;
power_data[2686] = 32'h00000086;
power_data[2687] = 32'h00000086;
power_data[2688] = 32'h00000086;
power_data[2689] = 32'h00000086;
power_data[2690] = 32'h00000086;
power_data[2691] = 32'h00000086;
power_data[2692] = 32'h00000086;
power_data[2693] = 32'h00000086;
power_data[2694] = 32'h00000086;
power_data[2695] = 32'h00000086;
power_data[2696] = 32'h00000086;
power_data[2697] = 32'h00000086;
power_data[2698] = 32'h00000086;
power_data[2699] = 32'h00000086;
power_data[2700] = 32'h00000086;
power_data[2701] = 32'h00000086;
power_data[2702] = 32'h00000086;
power_data[2703] = 32'h00000086;
power_data[2704] = 32'h00000086;
power_data[2705] = 32'h00000086;
power_data[2706] = 32'h00000086;
power_data[2707] = 32'h00000086;
power_data[2708] = 32'h00000086;
power_data[2709] = 32'h00000086;
power_data[2710] = 32'h00000086;
power_data[2711] = 32'h00000086;
power_data[2712] = 32'h00000086;
power_data[2713] = 32'h00000086;
power_data[2714] = 32'h00000086;
power_data[2715] = 32'h00000082;
power_data[2716] = 32'h00000069;
power_data[2717] = 32'h00000069;
power_data[2718] = 32'h00000069;
power_data[2719] = 32'h00000069;
power_data[2720] = 32'h00000069;
power_data[2721] = 32'h00000069;
power_data[2722] = 32'h00000069;
power_data[2723] = 32'h00000069;
power_data[2724] = 32'h00000069;
power_data[2725] = 32'h00000069;
power_data[2726] = 32'h00000069;
power_data[2727] = 32'h00000069;
power_data[2728] = 32'h00000069;
power_data[2729] = 32'h00000069;
power_data[2730] = 32'h00000069;
power_data[2731] = 32'h00000069;
power_data[2732] = 32'h00000069;
power_data[2733] = 32'h00000069;
power_data[2734] = 32'h00000069;
power_data[2735] = 32'h00000069;
power_data[2736] = 32'h00000069;
power_data[2737] = 32'h00000069;
power_data[2738] = 32'h00000069;
power_data[2739] = 32'h00000069;
power_data[2740] = 32'h00000069;
power_data[2741] = 32'h00000069;
power_data[2742] = 32'h00000069;
power_data[2743] = 32'h00000069;
power_data[2744] = 32'h00000069;
power_data[2745] = 32'h00000069;
power_data[2746] = 32'h00000069;
power_data[2747] = 32'h00000069;
power_data[2748] = 32'h00000069;
power_data[2749] = 32'h00000069;
power_data[2750] = 32'h00000069;
power_data[2751] = 32'h00000069;
power_data[2752] = 32'h00000069;
power_data[2753] = 32'h00000069;
power_data[2754] = 32'h00000069;
power_data[2755] = 32'h00000069;
power_data[2756] = 32'h00000069;
power_data[2757] = 32'h00000069;
power_data[2758] = 32'h00000069;
power_data[2759] = 32'h00000069;
power_data[2760] = 32'h00000069;
power_data[2761] = 32'h00000069;
power_data[2762] = 32'h00000069;
power_data[2763] = 32'h00000069;
power_data[2764] = 32'h00000069;
power_data[2765] = 32'h00000069;
power_data[2766] = 32'h00000069;
power_data[2767] = 32'h00000069;
power_data[2768] = 32'h00000069;
power_data[2769] = 32'h00000069;
power_data[2770] = 32'h00000069;
power_data[2771] = 32'h00000069;
power_data[2772] = 32'h00000069;
power_data[2773] = 32'h00000069;
power_data[2774] = 32'h00000069;
power_data[2775] = 32'h00000069;
power_data[2776] = 32'h00000069;
power_data[2777] = 32'h00000069;
power_data[2778] = 32'h00000069;
power_data[2779] = 32'h00000069;
power_data[2780] = 32'h00000069;
power_data[2781] = 32'h00000069;
power_data[2782] = 32'h00000069;
power_data[2783] = 32'h00000069;
power_data[2784] = 32'h00000069;
power_data[2785] = 32'h00000069;
power_data[2786] = 32'h0000077d;
power_data[2787] = 32'h00000942;
power_data[2788] = 32'h00000942;
power_data[2789] = 32'h00000942;
power_data[2790] = 32'h00000942;
power_data[2791] = 32'h00000942;
power_data[2792] = 32'h00000942;
power_data[2793] = 32'h00000942;
power_data[2794] = 32'h00000942;
power_data[2795] = 32'h00000942;
power_data[2796] = 32'h00000942;
power_data[2797] = 32'h00000942;
power_data[2798] = 32'h00000942;
power_data[2799] = 32'h00000942;
power_data[2800] = 32'h00000942;
power_data[2801] = 32'h00000942;
power_data[2802] = 32'h00000942;
power_data[2803] = 32'h00000942;
power_data[2804] = 32'h00000942;
power_data[2805] = 32'h00000942;
power_data[2806] = 32'h00000942;
power_data[2807] = 32'h00000942;
power_data[2808] = 32'h00000942;
power_data[2809] = 32'h00000942;
power_data[2810] = 32'h00000942;
power_data[2811] = 32'h00000942;
power_data[2812] = 32'h00000942;
power_data[2813] = 32'h00000942;
power_data[2814] = 32'h00000942;
power_data[2815] = 32'h00000232;
power_data[2816] = 32'h00000232;
power_data[2817] = 32'h00000232;
power_data[2818] = 32'h00000232;
power_data[2819] = 32'h00000232;
power_data[2820] = 32'h00000232;
power_data[2821] = 32'h00000232;
power_data[2822] = 32'h00000232;
power_data[2823] = 32'h00000232;
power_data[2824] = 32'h00000232;
power_data[2825] = 32'h00000232;
power_data[2826] = 32'h00000232;
power_data[2827] = 32'h00000232;
power_data[2828] = 32'h00000232;
power_data[2829] = 32'h00000232;
power_data[2830] = 32'h00000232;
power_data[2831] = 32'h00000232;
power_data[2832] = 32'h00000232;
power_data[2833] = 32'h00000232;
power_data[2834] = 32'h00000232;
power_data[2835] = 32'h00000232;
power_data[2836] = 32'h00000232;
power_data[2837] = 32'h00000232;
power_data[2838] = 32'h00000232;
power_data[2839] = 32'h00000232;
power_data[2840] = 32'h00000232;
power_data[2841] = 32'h00000232;
power_data[2842] = 32'h00000232;
power_data[2843] = 32'h00000232;
power_data[2844] = 32'h00000232;
power_data[2845] = 32'h00000232;
power_data[2846] = 32'h00000232;
power_data[2847] = 32'h00000232;
power_data[2848] = 32'h00000232;
power_data[2849] = 32'h00000232;
power_data[2850] = 32'h00000232;
power_data[2851] = 32'h00000232;
power_data[2852] = 32'h00000232;
power_data[2853] = 32'h00000232;
power_data[2854] = 32'h00000232;
power_data[2855] = 32'h00000232;
power_data[2856] = 32'h000013d3;
power_data[2857] = 32'h00002e41;
power_data[2858] = 32'h00002e41;
power_data[2859] = 32'h00002e41;
power_data[2860] = 32'h00002e41;
power_data[2861] = 32'h00002e41;
power_data[2862] = 32'h00002e41;
power_data[2863] = 32'h00002e41;
power_data[2864] = 32'h00002e41;
power_data[2865] = 32'h00002e41;
power_data[2866] = 32'h00002e41;
power_data[2867] = 32'h00002e41;
power_data[2868] = 32'h00002e41;
power_data[2869] = 32'h00002e41;
power_data[2870] = 32'h00002e41;
power_data[2871] = 32'h00002e41;
power_data[2872] = 32'h00002e41;
power_data[2873] = 32'h00002e41;
power_data[2874] = 32'h00002e41;
power_data[2875] = 32'h00002e41;
power_data[2876] = 32'h00002e41;
power_data[2877] = 32'h00002e41;
power_data[2878] = 32'h00002e41;
power_data[2879] = 32'h00002e41;
power_data[2880] = 32'h00002e41;
power_data[2881] = 32'h00002e41;
power_data[2882] = 32'h00002e41;
power_data[2883] = 32'h00002e41;
power_data[2884] = 32'h00002e41;
power_data[2885] = 32'h00002e41;
power_data[2886] = 32'h00002e41;
power_data[2887] = 32'h00002e41;
power_data[2888] = 32'h00002e41;
power_data[2889] = 32'h00002e41;
power_data[2890] = 32'h00002e41;
power_data[2891] = 32'h00002e41;
power_data[2892] = 32'h00002e41;
power_data[2893] = 32'h00002e41;
power_data[2894] = 32'h00002e41;
power_data[2895] = 32'h00002e41;
power_data[2896] = 32'h00002e41;
power_data[2897] = 32'h00002e41;
power_data[2898] = 32'h00002e41;
power_data[2899] = 32'h00002e41;
power_data[2900] = 32'h00002e41;
power_data[2901] = 32'h00002e41;
power_data[2902] = 32'h00002e41;
power_data[2903] = 32'h00002e41;
power_data[2904] = 32'h00002e41;
power_data[2905] = 32'h00002e41;
power_data[2906] = 32'h00002e41;
power_data[2907] = 32'h00002e41;
power_data[2908] = 32'h00002e41;
power_data[2909] = 32'h00002e41;
power_data[2910] = 32'h00002e41;
power_data[2911] = 32'h00002e41;
power_data[2912] = 32'h00002e41;
power_data[2913] = 32'h00002e41;
power_data[2914] = 32'h000009ab;
power_data[2915] = 32'h00000086;
power_data[2916] = 32'h00000086;
power_data[2917] = 32'h00000086;
power_data[2918] = 32'h00000086;
power_data[2919] = 32'h00000086;
power_data[2920] = 32'h00000086;
power_data[2921] = 32'h00000086;
power_data[2922] = 32'h00000086;
power_data[2923] = 32'h00000086;
power_data[2924] = 32'h00000086;
power_data[2925] = 32'h00000086;
power_data[2926] = 32'h00000086;
power_data[2927] = 32'h00000086;
power_data[2928] = 32'h00000086;
power_data[2929] = 32'h00000086;
power_data[2930] = 32'h00000086;
power_data[2931] = 32'h00000086;
power_data[2932] = 32'h00000086;
power_data[2933] = 32'h00000086;
power_data[2934] = 32'h00000086;
power_data[2935] = 32'h00000086;
power_data[2936] = 32'h00000086;
power_data[2937] = 32'h00000086;
power_data[2938] = 32'h00000086;
power_data[2939] = 32'h00000086;
power_data[2940] = 32'h00000086;
power_data[2941] = 32'h00000086;
power_data[2942] = 32'h00000086;
power_data[2943] = 32'h00000086;
power_data[2944] = 32'h00000086;
power_data[2945] = 32'h00000086;
power_data[2946] = 32'h00000086;
power_data[2947] = 32'h00000086;
power_data[2948] = 32'h00000086;
power_data[2949] = 32'h00000086;
power_data[2950] = 32'h00000086;
power_data[2951] = 32'h00000086;
power_data[2952] = 32'h00000086;
power_data[2953] = 32'h00000086;
power_data[2954] = 32'h00000086;
power_data[2955] = 32'h00000086;
power_data[2956] = 32'h00000086;
power_data[2957] = 32'h00000086;
power_data[2958] = 32'h00000086;
power_data[2959] = 32'h00000086;
power_data[2960] = 32'h00000086;
power_data[2961] = 32'h00000086;
power_data[2962] = 32'h00000086;
power_data[2963] = 32'h00000086;
power_data[2964] = 32'h00000086;
power_data[2965] = 32'h00000086;
power_data[2966] = 32'h00000086;
power_data[2967] = 32'h00000086;
power_data[2968] = 32'h00000086;
power_data[2969] = 32'h00000086;
power_data[2970] = 32'h00000086;
power_data[2971] = 32'h00000086;
power_data[2972] = 32'h00000086;
power_data[2973] = 32'h00000086;
power_data[2974] = 32'h00000086;
power_data[2975] = 32'h00000086;
power_data[2976] = 32'h00000086;
power_data[2977] = 32'h00000086;
power_data[2978] = 32'h00000086;
power_data[2979] = 32'h00000086;
power_data[2980] = 32'h00000086;
power_data[2981] = 32'h00000086;
power_data[2982] = 32'h00000086;
power_data[2983] = 32'h00000086;
power_data[2984] = 32'h00000086;
power_data[2985] = 32'h00000086;
power_data[2986] = 32'h00000086;
power_data[2987] = 32'h00000086;
power_data[2988] = 32'h00000086;
power_data[2989] = 32'h00000086;
power_data[2990] = 32'h00000086;
power_data[2991] = 32'h00000086;
power_data[2992] = 32'h00000086;
power_data[2993] = 32'h00000086;
power_data[2994] = 32'h00000086;
power_data[2995] = 32'h00000086;
power_data[2996] = 32'h00000086;
power_data[2997] = 32'h00000086;
power_data[2998] = 32'h00000086;
power_data[2999] = 32'h00000086;
power_data[3000] = 32'h00000086;
power_data[3001] = 32'h00000086;
power_data[3002] = 32'h00000086;
power_data[3003] = 32'h00000086;
power_data[3004] = 32'h00000086;
power_data[3005] = 32'h00000086;
power_data[3006] = 32'h00000086;
power_data[3007] = 32'h00000086;
power_data[3008] = 32'h00000086;
power_data[3009] = 32'h00000086;
power_data[3010] = 32'h00000086;
power_data[3011] = 32'h00000086;
power_data[3012] = 32'h00000086;
power_data[3013] = 32'h00000086;
power_data[3014] = 32'h00000086;
power_data[3015] = 32'h00000086;
power_data[3016] = 32'h00000086;
power_data[3017] = 32'h00000086;
power_data[3018] = 32'h00000086;
power_data[3019] = 32'h00000086;
power_data[3020] = 32'h00000086;
power_data[3021] = 32'h00000086;
power_data[3022] = 32'h00000086;
power_data[3023] = 32'h00000086;
power_data[3024] = 32'h00000086;
power_data[3025] = 32'h00000086;
power_data[3026] = 32'h00000086;
power_data[3027] = 32'h00000086;
power_data[3028] = 32'h00000086;
power_data[3029] = 32'h00000086;
power_data[3030] = 32'h00000086;
power_data[3031] = 32'h00000086;
power_data[3032] = 32'h00000086;
power_data[3033] = 32'h00000086;
power_data[3034] = 32'h00000086;
power_data[3035] = 32'h00000086;
power_data[3036] = 32'h00000086;
power_data[3037] = 32'h00000086;
power_data[3038] = 32'h00000086;
power_data[3039] = 32'h00000086;
power_data[3040] = 32'h00000086;
power_data[3041] = 32'h00000086;
power_data[3042] = 32'h00000086;
power_data[3043] = 32'h00000086;
power_data[3044] = 32'h00000086;
power_data[3045] = 32'h00000086;
power_data[3046] = 32'h00000086;
power_data[3047] = 32'h00000086;
power_data[3048] = 32'h00000086;
power_data[3049] = 32'h00000086;
power_data[3050] = 32'h00000086;
power_data[3051] = 32'h00000086;
power_data[3052] = 32'h00000086;
power_data[3053] = 32'h00000086;
power_data[3054] = 32'h00000086;
power_data[3055] = 32'h00000086;
power_data[3056] = 32'h00000086;
power_data[3057] = 32'h00000086;
power_data[3058] = 32'h00000086;
power_data[3059] = 32'h00000086;
power_data[3060] = 32'h00000086;
power_data[3061] = 32'h00000086;
power_data[3062] = 32'h00000086;
power_data[3063] = 32'h00000086;
power_data[3064] = 32'h00000086;
power_data[3065] = 32'h00000086;
power_data[3066] = 32'h00000086;
power_data[3067] = 32'h00000086;
power_data[3068] = 32'h00000086;
power_data[3069] = 32'h00000086;
power_data[3070] = 32'h00000086;
power_data[3071] = 32'h00000086;
power_data[3072] = 32'h00000086;
power_data[3073] = 32'h00000086;
power_data[3074] = 32'h00000086;
power_data[3075] = 32'h00000086;
power_data[3076] = 32'h00000086;
power_data[3077] = 32'h00000086;
power_data[3078] = 32'h00000086;
power_data[3079] = 32'h00000086;
power_data[3080] = 32'h00000086;
power_data[3081] = 32'h00000086;
power_data[3082] = 32'h00000086;
power_data[3083] = 32'h00000086;
power_data[3084] = 32'h00000086;
power_data[3085] = 32'h00000086;
power_data[3086] = 32'h00000086;
power_data[3087] = 32'h00000086;
power_data[3088] = 32'h00000086;
power_data[3089] = 32'h00000086;
power_data[3090] = 32'h00000086;
power_data[3091] = 32'h00000086;
power_data[3092] = 32'h00000086;
power_data[3093] = 32'h00000086;
power_data[3094] = 32'h00000086;
power_data[3095] = 32'h00000086;
power_data[3096] = 32'h00000086;
power_data[3097] = 32'h00000086;
power_data[3098] = 32'h00000086;
power_data[3099] = 32'h00000086;
power_data[3100] = 32'h00000086;
power_data[3101] = 32'h00000086;
power_data[3102] = 32'h00000086;
power_data[3103] = 32'h00000086;
power_data[3104] = 32'h00000086;
power_data[3105] = 32'h00000086;
power_data[3106] = 32'h00000086;
power_data[3107] = 32'h00000086;
power_data[3108] = 32'h00000086;
power_data[3109] = 32'h00000086;
power_data[3110] = 32'h00000086;
power_data[3111] = 32'h00000086;
power_data[3112] = 32'h00000086;
power_data[3113] = 32'h00000086;
power_data[3114] = 32'h00000086;
power_data[3115] = 32'h00000086;
power_data[3116] = 32'h00000086;
power_data[3117] = 32'h00000086;
power_data[3118] = 32'h00000086;
power_data[3119] = 32'h00000086;
power_data[3120] = 32'h00000086;
power_data[3121] = 32'h00000086;
power_data[3122] = 32'h00000086;
power_data[3123] = 32'h00000086;
power_data[3124] = 32'h00000086;
power_data[3125] = 32'h00000086;
power_data[3126] = 32'h00000086;
power_data[3127] = 32'h00000086;
power_data[3128] = 32'h00000086;
power_data[3129] = 32'h00000086;
power_data[3130] = 32'h00000086;
power_data[3131] = 32'h00000086;
power_data[3132] = 32'h00000086;
power_data[3133] = 32'h00000086;
power_data[3134] = 32'h00000086;
power_data[3135] = 32'h00000086;
power_data[3136] = 32'h00000086;
power_data[3137] = 32'h00000086;
power_data[3138] = 32'h00000086;
power_data[3139] = 32'h00000086;
power_data[3140] = 32'h00000086;
power_data[3141] = 32'h00000086;
power_data[3142] = 32'h00000086;
power_data[3143] = 32'h00000086;
power_data[3144] = 32'h00000086;
power_data[3145] = 32'h00000086;
power_data[3146] = 32'h00000086;
power_data[3147] = 32'h00000086;
power_data[3148] = 32'h00000086;
power_data[3149] = 32'h00000086;
power_data[3150] = 32'h00000086;
power_data[3151] = 32'h00000086;
power_data[3152] = 32'h00000086;
power_data[3153] = 32'h00000086;
power_data[3154] = 32'h00000086;
power_data[3155] = 32'h00000086;
power_data[3156] = 32'h00000086;
power_data[3157] = 32'h00000086;
power_data[3158] = 32'h00000086;
power_data[3159] = 32'h00000086;
power_data[3160] = 32'h00000086;
power_data[3161] = 32'h00000086;
power_data[3162] = 32'h00000086;
power_data[3163] = 32'h00000086;
power_data[3164] = 32'h00000086;
power_data[3165] = 32'h00000086;
power_data[3166] = 32'h00000086;
power_data[3167] = 32'h00000086;
power_data[3168] = 32'h00000086;
power_data[3169] = 32'h00000086;
power_data[3170] = 32'h00000086;
power_data[3171] = 32'h00000086;
power_data[3172] = 32'h00000086;
power_data[3173] = 32'h00000086;
power_data[3174] = 32'h00000086;
power_data[3175] = 32'h00000086;
power_data[3176] = 32'h00000086;
power_data[3177] = 32'h00000086;
power_data[3178] = 32'h00000086;
power_data[3179] = 32'h00000086;
power_data[3180] = 32'h00000086;
power_data[3181] = 32'h00000086;
power_data[3182] = 32'h00000086;
power_data[3183] = 32'h00000086;
power_data[3184] = 32'h00000086;
power_data[3185] = 32'h00000086;
power_data[3186] = 32'h00000086;
power_data[3187] = 32'h00000086;
power_data[3188] = 32'h00000086;
power_data[3189] = 32'h00000086;
power_data[3190] = 32'h00000086;
power_data[3191] = 32'h00000086;
power_data[3192] = 32'h00000086;
power_data[3193] = 32'h00000086;
power_data[3194] = 32'h00000086;
power_data[3195] = 32'h00000086;
power_data[3196] = 32'h00000086;
power_data[3197] = 32'h00000086;
power_data[3198] = 32'h00000086;
power_data[3199] = 32'h00000086;
power_data[3200] = 32'h00000086;
power_data[3201] = 32'h00000086;
power_data[3202] = 32'h00000086;
power_data[3203] = 32'h00000086;
power_data[3204] = 32'h00000086;
power_data[3205] = 32'h00000086;
power_data[3206] = 32'h00000086;
power_data[3207] = 32'h00000086;
power_data[3208] = 32'h00000086;
power_data[3209] = 32'h00000086;
power_data[3210] = 32'h00000086;
power_data[3211] = 32'h00000086;
power_data[3212] = 32'h00000086;
power_data[3213] = 32'h00000086;
power_data[3214] = 32'h00000086;
power_data[3215] = 32'h00000086;
power_data[3216] = 32'h00000086;
power_data[3217] = 32'h00000086;
power_data[3218] = 32'h00000086;
power_data[3219] = 32'h00000086;
power_data[3220] = 32'h00000086;
power_data[3221] = 32'h00000086;
power_data[3222] = 32'h00000086;
power_data[3223] = 32'h00000086;
power_data[3224] = 32'h00000086;
power_data[3225] = 32'h00000086;
power_data[3226] = 32'h00000086;
power_data[3227] = 32'h00000082;
power_data[3228] = 32'h00000069;
power_data[3229] = 32'h00000069;
power_data[3230] = 32'h00000069;
power_data[3231] = 32'h00000069;
power_data[3232] = 32'h00000069;
power_data[3233] = 32'h00000069;
power_data[3234] = 32'h00000069;
power_data[3235] = 32'h00000069;
power_data[3236] = 32'h00000069;
power_data[3237] = 32'h00000069;
power_data[3238] = 32'h00000069;
power_data[3239] = 32'h00000069;
power_data[3240] = 32'h00000069;
power_data[3241] = 32'h00000069;
power_data[3242] = 32'h00000069;
power_data[3243] = 32'h00000069;
power_data[3244] = 32'h00000069;
power_data[3245] = 32'h00000069;
power_data[3246] = 32'h00000069;
power_data[3247] = 32'h00000069;
power_data[3248] = 32'h00000069;
power_data[3249] = 32'h00000069;
power_data[3250] = 32'h00000069;
power_data[3251] = 32'h00000069;
power_data[3252] = 32'h00000069;
power_data[3253] = 32'h00000069;
power_data[3254] = 32'h00000069;
power_data[3255] = 32'h00000069;
power_data[3256] = 32'h00000069;
power_data[3257] = 32'h00000069;
power_data[3258] = 32'h00000069;
power_data[3259] = 32'h00000069;
power_data[3260] = 32'h00000069;
power_data[3261] = 32'h00000069;
power_data[3262] = 32'h00000069;
power_data[3263] = 32'h00000069;
power_data[3264] = 32'h00000069;
power_data[3265] = 32'h00000069;
power_data[3266] = 32'h00000069;
power_data[3267] = 32'h00000069;
power_data[3268] = 32'h00000069;
power_data[3269] = 32'h00000069;
power_data[3270] = 32'h00000069;
power_data[3271] = 32'h00000069;
power_data[3272] = 32'h00000069;
power_data[3273] = 32'h00000069;
power_data[3274] = 32'h00000069;
power_data[3275] = 32'h00000069;
power_data[3276] = 32'h00000069;
power_data[3277] = 32'h00000069;
power_data[3278] = 32'h00000069;
power_data[3279] = 32'h00000069;
power_data[3280] = 32'h00000069;
power_data[3281] = 32'h00000069;
power_data[3282] = 32'h00000069;
power_data[3283] = 32'h00000069;
power_data[3284] = 32'h00000069;
power_data[3285] = 32'h00000069;
power_data[3286] = 32'h00000069;
power_data[3287] = 32'h00000069;
power_data[3288] = 32'h00000069;
power_data[3289] = 32'h00000069;
power_data[3290] = 32'h00000069;
power_data[3291] = 32'h00000069;
power_data[3292] = 32'h00000069;
power_data[3293] = 32'h00000069;
power_data[3294] = 32'h00000069;
power_data[3295] = 32'h00000069;
power_data[3296] = 32'h00000069;
power_data[3297] = 32'h00000069;
power_data[3298] = 32'h0000077d;
power_data[3299] = 32'h00000942;
power_data[3300] = 32'h00000942;
power_data[3301] = 32'h00000942;
power_data[3302] = 32'h00000942;
power_data[3303] = 32'h00000942;
power_data[3304] = 32'h00000942;
power_data[3305] = 32'h00000942;
power_data[3306] = 32'h00000942;
power_data[3307] = 32'h00000942;
power_data[3308] = 32'h00000942;
power_data[3309] = 32'h00000942;
power_data[3310] = 32'h00000942;
power_data[3311] = 32'h00000942;
power_data[3312] = 32'h00000942;
power_data[3313] = 32'h00000942;
power_data[3314] = 32'h00000942;
power_data[3315] = 32'h00000942;
power_data[3316] = 32'h00000942;
power_data[3317] = 32'h00000942;
power_data[3318] = 32'h00000942;
power_data[3319] = 32'h00000942;
power_data[3320] = 32'h00000942;
power_data[3321] = 32'h00000942;
power_data[3322] = 32'h00000942;
power_data[3323] = 32'h00000942;
power_data[3324] = 32'h00000942;
power_data[3325] = 32'h00000942;
power_data[3326] = 32'h00000942;
power_data[3327] = 32'h00000232;
power_data[3328] = 32'h00000232;
power_data[3329] = 32'h00000232;
power_data[3330] = 32'h00000232;
power_data[3331] = 32'h00000232;
power_data[3332] = 32'h00000232;
power_data[3333] = 32'h00000232;
power_data[3334] = 32'h00000232;
power_data[3335] = 32'h00000232;
power_data[3336] = 32'h00000232;
power_data[3337] = 32'h00000232;
power_data[3338] = 32'h00000232;
power_data[3339] = 32'h00000232;
power_data[3340] = 32'h00000232;
power_data[3341] = 32'h00000232;
power_data[3342] = 32'h00000232;
power_data[3343] = 32'h00000232;
power_data[3344] = 32'h00000232;
power_data[3345] = 32'h00000232;
power_data[3346] = 32'h00000232;
power_data[3347] = 32'h00000232;
power_data[3348] = 32'h00000232;
power_data[3349] = 32'h00000232;
power_data[3350] = 32'h00000232;
power_data[3351] = 32'h00000232;
power_data[3352] = 32'h00000232;
power_data[3353] = 32'h00000232;
power_data[3354] = 32'h00000232;
power_data[3355] = 32'h00000232;
power_data[3356] = 32'h00000232;
power_data[3357] = 32'h00000232;
power_data[3358] = 32'h00000232;
power_data[3359] = 32'h00000232;
power_data[3360] = 32'h00000232;
power_data[3361] = 32'h00000232;
power_data[3362] = 32'h00000232;
power_data[3363] = 32'h00000232;
power_data[3364] = 32'h00000232;
power_data[3365] = 32'h00000232;
power_data[3366] = 32'h00000232;
power_data[3367] = 32'h00000232;
power_data[3368] = 32'h000013d3;
power_data[3369] = 32'h00002e41;
power_data[3370] = 32'h00002e41;
power_data[3371] = 32'h00002e41;
power_data[3372] = 32'h00002e41;
power_data[3373] = 32'h00002e41;
power_data[3374] = 32'h00002e41;
power_data[3375] = 32'h00002e41;
power_data[3376] = 32'h00002e41;
power_data[3377] = 32'h00002e41;
power_data[3378] = 32'h00002e41;
power_data[3379] = 32'h00002e41;
power_data[3380] = 32'h00002e41;
power_data[3381] = 32'h00002e41;
power_data[3382] = 32'h00002e41;
power_data[3383] = 32'h00002e41;
power_data[3384] = 32'h00002e41;
power_data[3385] = 32'h00002e41;
power_data[3386] = 32'h00002e41;
power_data[3387] = 32'h00002e41;
power_data[3388] = 32'h00002e41;
power_data[3389] = 32'h00002e41;
power_data[3390] = 32'h00002e41;
power_data[3391] = 32'h00002e41;
power_data[3392] = 32'h00002e41;
power_data[3393] = 32'h00002e41;
power_data[3394] = 32'h00002e41;
power_data[3395] = 32'h00002e41;
power_data[3396] = 32'h00002e41;
power_data[3397] = 32'h00002e41;
power_data[3398] = 32'h00002e41;
power_data[3399] = 32'h00002e41;
power_data[3400] = 32'h00002e41;
power_data[3401] = 32'h00002e41;
power_data[3402] = 32'h00002e41;
power_data[3403] = 32'h00002e41;
power_data[3404] = 32'h00002e41;
power_data[3405] = 32'h00002e41;
power_data[3406] = 32'h00002e41;
power_data[3407] = 32'h00002e41;
power_data[3408] = 32'h00002e41;
power_data[3409] = 32'h00002e41;
power_data[3410] = 32'h00002e41;
power_data[3411] = 32'h00002e41;
power_data[3412] = 32'h00002e41;
power_data[3413] = 32'h00002e41;
power_data[3414] = 32'h00002e41;
power_data[3415] = 32'h00002e41;
power_data[3416] = 32'h00002e41;
power_data[3417] = 32'h00002e41;
power_data[3418] = 32'h00002e41;
power_data[3419] = 32'h00002e41;
power_data[3420] = 32'h00002e41;
power_data[3421] = 32'h00002e41;
power_data[3422] = 32'h00002e41;
power_data[3423] = 32'h00002e41;
power_data[3424] = 32'h00002e41;
power_data[3425] = 32'h00002e41;
power_data[3426] = 32'h000009ab;
power_data[3427] = 32'h00000086;
power_data[3428] = 32'h00000086;
power_data[3429] = 32'h00000086;
power_data[3430] = 32'h00000086;
power_data[3431] = 32'h00000086;
power_data[3432] = 32'h00000086;
power_data[3433] = 32'h00000086;
power_data[3434] = 32'h00000086;
power_data[3435] = 32'h00000086;
power_data[3436] = 32'h00000086;
power_data[3437] = 32'h00000086;
power_data[3438] = 32'h00000086;
power_data[3439] = 32'h00000086;
power_data[3440] = 32'h00000086;
power_data[3441] = 32'h00000086;
power_data[3442] = 32'h00000086;
power_data[3443] = 32'h00000086;
power_data[3444] = 32'h00000086;
power_data[3445] = 32'h00000086;
power_data[3446] = 32'h00000086;
power_data[3447] = 32'h00000086;
power_data[3448] = 32'h00000086;
power_data[3449] = 32'h00000086;
power_data[3450] = 32'h00000086;
power_data[3451] = 32'h00000086;
power_data[3452] = 32'h00000086;
power_data[3453] = 32'h00000086;
power_data[3454] = 32'h00000086;
power_data[3455] = 32'h00000086;
power_data[3456] = 32'h00000086;
power_data[3457] = 32'h00000086;
power_data[3458] = 32'h00000086;
power_data[3459] = 32'h00000086;
power_data[3460] = 32'h00000086;
power_data[3461] = 32'h00000086;
power_data[3462] = 32'h00000086;
power_data[3463] = 32'h00000086;
power_data[3464] = 32'h00000086;
power_data[3465] = 32'h00000086;
power_data[3466] = 32'h00000086;
power_data[3467] = 32'h00000086;
power_data[3468] = 32'h00000086;
power_data[3469] = 32'h00000086;
power_data[3470] = 32'h00000086;
power_data[3471] = 32'h00000086;
power_data[3472] = 32'h00000086;
power_data[3473] = 32'h00000086;
power_data[3474] = 32'h00000086;
power_data[3475] = 32'h00000086;
power_data[3476] = 32'h00000086;
power_data[3477] = 32'h00000086;
power_data[3478] = 32'h00000086;
power_data[3479] = 32'h00000086;
power_data[3480] = 32'h00000086;
power_data[3481] = 32'h00000086;
power_data[3482] = 32'h00000086;
power_data[3483] = 32'h00000086;
power_data[3484] = 32'h00000086;
power_data[3485] = 32'h00000086;
power_data[3486] = 32'h00000086;
power_data[3487] = 32'h00000086;
power_data[3488] = 32'h00000086;
power_data[3489] = 32'h00000086;
power_data[3490] = 32'h00000086;
power_data[3491] = 32'h00000086;
power_data[3492] = 32'h00000086;
power_data[3493] = 32'h00000086;
power_data[3494] = 32'h00000086;
power_data[3495] = 32'h00000086;
power_data[3496] = 32'h00000086;
power_data[3497] = 32'h00000086;
power_data[3498] = 32'h00000086;
power_data[3499] = 32'h00000086;
power_data[3500] = 32'h00000086;
power_data[3501] = 32'h00000086;
power_data[3502] = 32'h00000086;
power_data[3503] = 32'h00000086;
power_data[3504] = 32'h00000086;
power_data[3505] = 32'h00000086;
power_data[3506] = 32'h00000086;
power_data[3507] = 32'h00000086;
power_data[3508] = 32'h00000086;
power_data[3509] = 32'h00000086;
power_data[3510] = 32'h00000086;
power_data[3511] = 32'h00000086;
power_data[3512] = 32'h00000086;
power_data[3513] = 32'h00000086;
power_data[3514] = 32'h00000086;
power_data[3515] = 32'h00000086;
power_data[3516] = 32'h00000086;
power_data[3517] = 32'h00000086;
power_data[3518] = 32'h00000086;
power_data[3519] = 32'h00000086;
power_data[3520] = 32'h00000086;
power_data[3521] = 32'h00000086;
power_data[3522] = 32'h00000086;
power_data[3523] = 32'h00000086;
power_data[3524] = 32'h00000086;
power_data[3525] = 32'h00000086;
power_data[3526] = 32'h00000086;
power_data[3527] = 32'h00000086;
power_data[3528] = 32'h00000086;
power_data[3529] = 32'h00000086;
power_data[3530] = 32'h00000086;
power_data[3531] = 32'h00000086;
power_data[3532] = 32'h00000086;
power_data[3533] = 32'h00000086;
power_data[3534] = 32'h00000086;
power_data[3535] = 32'h00000086;
power_data[3536] = 32'h00000086;
power_data[3537] = 32'h00000086;
power_data[3538] = 32'h00000086;
power_data[3539] = 32'h00000086;
power_data[3540] = 32'h00000086;
power_data[3541] = 32'h00000086;
power_data[3542] = 32'h00000086;
power_data[3543] = 32'h00000086;
power_data[3544] = 32'h00000086;
power_data[3545] = 32'h00000086;
power_data[3546] = 32'h00000086;
power_data[3547] = 32'h00000086;
power_data[3548] = 32'h00000086;
power_data[3549] = 32'h00000086;
power_data[3550] = 32'h00000086;
power_data[3551] = 32'h00000086;
power_data[3552] = 32'h00000086;
power_data[3553] = 32'h00000086;
power_data[3554] = 32'h00000086;
power_data[3555] = 32'h00000086;
power_data[3556] = 32'h00000086;
power_data[3557] = 32'h00000086;
power_data[3558] = 32'h00000086;
power_data[3559] = 32'h00000086;
power_data[3560] = 32'h00000086;
power_data[3561] = 32'h00000086;
power_data[3562] = 32'h00000086;
power_data[3563] = 32'h00000086;
power_data[3564] = 32'h00000086;
power_data[3565] = 32'h00000086;
power_data[3566] = 32'h00000086;
power_data[3567] = 32'h00000086;
power_data[3568] = 32'h00000086;
power_data[3569] = 32'h00000086;
power_data[3570] = 32'h00000086;
power_data[3571] = 32'h00000086;
power_data[3572] = 32'h00000086;
power_data[3573] = 32'h00000086;
power_data[3574] = 32'h00000086;
power_data[3575] = 32'h00000086;
power_data[3576] = 32'h00000086;
power_data[3577] = 32'h00000086;
power_data[3578] = 32'h00000086;
power_data[3579] = 32'h00000086;
power_data[3580] = 32'h00000086;
power_data[3581] = 32'h00000086;
power_data[3582] = 32'h00000086;
power_data[3583] = 32'h00000086;
power_data[3584] = 32'h00000086;
power_data[3585] = 32'h00000086;
power_data[3586] = 32'h00000086;
power_data[3587] = 32'h00000086;
power_data[3588] = 32'h00000086;
power_data[3589] = 32'h00000086;
power_data[3590] = 32'h00000086;
power_data[3591] = 32'h00000086;
power_data[3592] = 32'h00000086;
power_data[3593] = 32'h00000086;
power_data[3594] = 32'h00000086;
power_data[3595] = 32'h00000086;
power_data[3596] = 32'h00000086;
power_data[3597] = 32'h00000086;
power_data[3598] = 32'h00000086;
power_data[3599] = 32'h00000086;
power_data[3600] = 32'h00000086;
power_data[3601] = 32'h00000086;
power_data[3602] = 32'h00000086;
power_data[3603] = 32'h00000086;
power_data[3604] = 32'h00000086;
power_data[3605] = 32'h00000086;
power_data[3606] = 32'h00000086;
power_data[3607] = 32'h00000086;
power_data[3608] = 32'h00000086;
power_data[3609] = 32'h00000086;
power_data[3610] = 32'h00000086;
power_data[3611] = 32'h00000086;
power_data[3612] = 32'h00000086;
power_data[3613] = 32'h00000086;
power_data[3614] = 32'h00000086;
power_data[3615] = 32'h00000086;
power_data[3616] = 32'h00000086;
power_data[3617] = 32'h00000086;
power_data[3618] = 32'h00000086;
power_data[3619] = 32'h00000086;
power_data[3620] = 32'h00000086;
power_data[3621] = 32'h00000086;
power_data[3622] = 32'h00000086;
power_data[3623] = 32'h00000086;
power_data[3624] = 32'h00000086;
power_data[3625] = 32'h00000086;
power_data[3626] = 32'h00000086;
power_data[3627] = 32'h00000086;
power_data[3628] = 32'h00000086;
power_data[3629] = 32'h00000086;
power_data[3630] = 32'h00000086;
power_data[3631] = 32'h00000086;
power_data[3632] = 32'h00000086;
power_data[3633] = 32'h00000086;
power_data[3634] = 32'h00000086;
power_data[3635] = 32'h00000086;
power_data[3636] = 32'h00000086;
power_data[3637] = 32'h00000086;
power_data[3638] = 32'h00000086;
power_data[3639] = 32'h00000086;
power_data[3640] = 32'h00000086;
power_data[3641] = 32'h00000086;
power_data[3642] = 32'h00000086;
power_data[3643] = 32'h00000086;
power_data[3644] = 32'h00000086;
power_data[3645] = 32'h00000086;
power_data[3646] = 32'h00000086;
power_data[3647] = 32'h00000086;
power_data[3648] = 32'h00000086;
power_data[3649] = 32'h00000086;
power_data[3650] = 32'h00000086;
power_data[3651] = 32'h00000086;
power_data[3652] = 32'h00000086;
power_data[3653] = 32'h00000086;
power_data[3654] = 32'h00000086;
power_data[3655] = 32'h00000086;
power_data[3656] = 32'h00000086;
power_data[3657] = 32'h00000086;
power_data[3658] = 32'h00000086;
power_data[3659] = 32'h00000086;
power_data[3660] = 32'h00000086;
power_data[3661] = 32'h00000086;
power_data[3662] = 32'h00000086;
power_data[3663] = 32'h00000086;
power_data[3664] = 32'h00000086;
power_data[3665] = 32'h00000086;
power_data[3666] = 32'h00000086;
power_data[3667] = 32'h00000086;
power_data[3668] = 32'h00000086;
power_data[3669] = 32'h00000086;
power_data[3670] = 32'h00000086;
power_data[3671] = 32'h00000086;
power_data[3672] = 32'h00000086;
power_data[3673] = 32'h00000086;
power_data[3674] = 32'h00000086;
power_data[3675] = 32'h00000086;
power_data[3676] = 32'h00000086;
power_data[3677] = 32'h00000086;
power_data[3678] = 32'h00000086;
power_data[3679] = 32'h00000086;
power_data[3680] = 32'h00000086;
power_data[3681] = 32'h00000086;
power_data[3682] = 32'h00000086;
power_data[3683] = 32'h00000086;
power_data[3684] = 32'h00000086;
power_data[3685] = 32'h00000086;
power_data[3686] = 32'h00000086;
power_data[3687] = 32'h00000086;
power_data[3688] = 32'h00000086;
power_data[3689] = 32'h00000086;
power_data[3690] = 32'h00000086;
power_data[3691] = 32'h00000086;
power_data[3692] = 32'h00000086;
power_data[3693] = 32'h00000086;
power_data[3694] = 32'h00000086;
power_data[3695] = 32'h00000086;
power_data[3696] = 32'h00000086;
power_data[3697] = 32'h00000086;
power_data[3698] = 32'h00000086;
power_data[3699] = 32'h00000086;
power_data[3700] = 32'h00000086;
power_data[3701] = 32'h00000086;
power_data[3702] = 32'h00000086;
power_data[3703] = 32'h00000086;
power_data[3704] = 32'h00000086;
power_data[3705] = 32'h00000086;
power_data[3706] = 32'h00000086;
power_data[3707] = 32'h00000086;
power_data[3708] = 32'h00000086;
power_data[3709] = 32'h00000086;
power_data[3710] = 32'h00000086;
power_data[3711] = 32'h00000086;
power_data[3712] = 32'h00000086;
power_data[3713] = 32'h00000086;
power_data[3714] = 32'h00000086;
power_data[3715] = 32'h00000086;
power_data[3716] = 32'h00000086;
power_data[3717] = 32'h00000086;
power_data[3718] = 32'h00000086;
power_data[3719] = 32'h00000086;
power_data[3720] = 32'h00000086;
power_data[3721] = 32'h00000086;
power_data[3722] = 32'h00000086;
power_data[3723] = 32'h00000086;
power_data[3724] = 32'h00000086;
power_data[3725] = 32'h00000086;
power_data[3726] = 32'h00000086;
power_data[3727] = 32'h00000086;
power_data[3728] = 32'h00000086;
power_data[3729] = 32'h00000086;
power_data[3730] = 32'h00000086;
power_data[3731] = 32'h00000086;
power_data[3732] = 32'h00000086;
power_data[3733] = 32'h00000086;
power_data[3734] = 32'h00000086;
power_data[3735] = 32'h00000086;
power_data[3736] = 32'h00000086;
power_data[3737] = 32'h00000086;
power_data[3738] = 32'h00000086;
power_data[3739] = 32'h00000082;
power_data[3740] = 32'h00000069;
power_data[3741] = 32'h00000069;
power_data[3742] = 32'h00000069;
power_data[3743] = 32'h00000069;
power_data[3744] = 32'h00000069;
power_data[3745] = 32'h00000069;
power_data[3746] = 32'h00000069;
power_data[3747] = 32'h00000069;
power_data[3748] = 32'h00000069;
power_data[3749] = 32'h00000069;
power_data[3750] = 32'h00000069;
power_data[3751] = 32'h00000069;
power_data[3752] = 32'h00000069;
power_data[3753] = 32'h00000069;
power_data[3754] = 32'h00000069;
power_data[3755] = 32'h00000069;
power_data[3756] = 32'h00000069;
power_data[3757] = 32'h00000069;
power_data[3758] = 32'h00000069;
power_data[3759] = 32'h00000069;
power_data[3760] = 32'h00000069;
power_data[3761] = 32'h00000069;
power_data[3762] = 32'h00000069;
power_data[3763] = 32'h00000069;
power_data[3764] = 32'h00000069;
power_data[3765] = 32'h00000069;
power_data[3766] = 32'h00000069;
power_data[3767] = 32'h00000069;
power_data[3768] = 32'h00000069;
power_data[3769] = 32'h00000069;
power_data[3770] = 32'h00000069;
power_data[3771] = 32'h00000069;
power_data[3772] = 32'h00000069;
power_data[3773] = 32'h00000069;
power_data[3774] = 32'h00000069;
power_data[3775] = 32'h00000069;
power_data[3776] = 32'h00000069;
power_data[3777] = 32'h00000069;
power_data[3778] = 32'h00000069;
power_data[3779] = 32'h00000069;
power_data[3780] = 32'h00000069;
power_data[3781] = 32'h00000069;
power_data[3782] = 32'h00000069;
power_data[3783] = 32'h00000069;
power_data[3784] = 32'h00000069;
power_data[3785] = 32'h00000069;
power_data[3786] = 32'h00000069;
power_data[3787] = 32'h00000069;
power_data[3788] = 32'h00000069;
power_data[3789] = 32'h00000069;
power_data[3790] = 32'h00000069;
power_data[3791] = 32'h00000069;
power_data[3792] = 32'h00000069;
power_data[3793] = 32'h00000069;
power_data[3794] = 32'h00000069;
power_data[3795] = 32'h00000069;
power_data[3796] = 32'h00000069;
power_data[3797] = 32'h00000069;
power_data[3798] = 32'h00000069;
power_data[3799] = 32'h00000069;
power_data[3800] = 32'h00000069;
power_data[3801] = 32'h00000069;
power_data[3802] = 32'h00000069;
power_data[3803] = 32'h00000069;
power_data[3804] = 32'h00000069;
power_data[3805] = 32'h00000069;
power_data[3806] = 32'h00000069;
power_data[3807] = 32'h00000069;
power_data[3808] = 32'h00000069;
power_data[3809] = 32'h00000069;
power_data[3810] = 32'h0000077d;
power_data[3811] = 32'h00000942;
power_data[3812] = 32'h00000942;
power_data[3813] = 32'h00000942;
power_data[3814] = 32'h00000942;
power_data[3815] = 32'h00000942;
power_data[3816] = 32'h00000942;
power_data[3817] = 32'h00000942;
power_data[3818] = 32'h00000942;
power_data[3819] = 32'h00000942;
power_data[3820] = 32'h00000942;
power_data[3821] = 32'h00000942;
power_data[3822] = 32'h00000942;
power_data[3823] = 32'h00000942;
power_data[3824] = 32'h00000942;
power_data[3825] = 32'h00000942;
power_data[3826] = 32'h00000942;
power_data[3827] = 32'h00000942;
power_data[3828] = 32'h00000942;
power_data[3829] = 32'h00000942;
power_data[3830] = 32'h00000942;
power_data[3831] = 32'h00000942;
power_data[3832] = 32'h00000942;
power_data[3833] = 32'h00000942;
power_data[3834] = 32'h00000942;
power_data[3835] = 32'h00000942;
power_data[3836] = 32'h00000942;
power_data[3837] = 32'h00000942;
power_data[3838] = 32'h00000942;
power_data[3839] = 32'h00000232;
power_data[3840] = 32'h00000232;
power_data[3841] = 32'h00000232;
power_data[3842] = 32'h00000232;
power_data[3843] = 32'h00000232;
power_data[3844] = 32'h00000232;
power_data[3845] = 32'h00000232;
power_data[3846] = 32'h00000232;
power_data[3847] = 32'h00000232;
power_data[3848] = 32'h00000232;
power_data[3849] = 32'h00000232;
power_data[3850] = 32'h00000232;
power_data[3851] = 32'h00000232;
power_data[3852] = 32'h00000232;
power_data[3853] = 32'h00000232;
power_data[3854] = 32'h00000232;
power_data[3855] = 32'h00000232;
power_data[3856] = 32'h00000232;
power_data[3857] = 32'h00000232;
power_data[3858] = 32'h00000232;
power_data[3859] = 32'h00000232;
power_data[3860] = 32'h00000232;
power_data[3861] = 32'h00000232;
power_data[3862] = 32'h00000232;
power_data[3863] = 32'h00000232;
power_data[3864] = 32'h00000232;
power_data[3865] = 32'h00000232;
power_data[3866] = 32'h00000232;
power_data[3867] = 32'h00000232;
power_data[3868] = 32'h00000232;
power_data[3869] = 32'h00000232;
power_data[3870] = 32'h00000232;
power_data[3871] = 32'h00000232;
power_data[3872] = 32'h00000232;
power_data[3873] = 32'h00000232;
power_data[3874] = 32'h00000232;
power_data[3875] = 32'h00000232;
power_data[3876] = 32'h00000232;
power_data[3877] = 32'h00000232;
power_data[3878] = 32'h00000232;
power_data[3879] = 32'h00000232;
power_data[3880] = 32'h000013d3;
power_data[3881] = 32'h00002e41;
power_data[3882] = 32'h00002e41;
power_data[3883] = 32'h00002e41;
power_data[3884] = 32'h00002e41;
power_data[3885] = 32'h00002e41;
power_data[3886] = 32'h00002e41;
power_data[3887] = 32'h00002e41;
power_data[3888] = 32'h00002e41;
power_data[3889] = 32'h00002e41;
power_data[3890] = 32'h00002e41;
power_data[3891] = 32'h00002e41;
power_data[3892] = 32'h00002e41;
power_data[3893] = 32'h00002e41;
power_data[3894] = 32'h00002e41;
power_data[3895] = 32'h00002e41;
power_data[3896] = 32'h00002e41;
power_data[3897] = 32'h00002e41;
power_data[3898] = 32'h00002e41;
power_data[3899] = 32'h00002e41;
power_data[3900] = 32'h00002e41;
power_data[3901] = 32'h00002e41;
power_data[3902] = 32'h00002e41;
power_data[3903] = 32'h00002e41;
power_data[3904] = 32'h00002e41;
power_data[3905] = 32'h00002e41;
power_data[3906] = 32'h00002e41;
power_data[3907] = 32'h00002e41;
power_data[3908] = 32'h00002e41;
power_data[3909] = 32'h00002e41;
power_data[3910] = 32'h00002e41;
power_data[3911] = 32'h00002e41;
power_data[3912] = 32'h00002e41;
power_data[3913] = 32'h00002e41;
power_data[3914] = 32'h00002e41;
power_data[3915] = 32'h00002e41;
power_data[3916] = 32'h00002e41;
power_data[3917] = 32'h00002e41;
power_data[3918] = 32'h00002e41;
power_data[3919] = 32'h00002e41;
power_data[3920] = 32'h00002e41;
power_data[3921] = 32'h00002e41;
power_data[3922] = 32'h00002e41;
power_data[3923] = 32'h00002e41;
power_data[3924] = 32'h00002e41;
power_data[3925] = 32'h00002e41;
power_data[3926] = 32'h00002e41;
power_data[3927] = 32'h00002e41;
power_data[3928] = 32'h00002e41;
power_data[3929] = 32'h00002e41;
power_data[3930] = 32'h00002e41;
power_data[3931] = 32'h00002e41;
power_data[3932] = 32'h00002e41;
power_data[3933] = 32'h00002e41;
power_data[3934] = 32'h00002e41;
power_data[3935] = 32'h00002e41;
power_data[3936] = 32'h00002e41;
power_data[3937] = 32'h00002e41;
power_data[3938] = 32'h000009ab;
power_data[3939] = 32'h00000086;
power_data[3940] = 32'h00000086;
power_data[3941] = 32'h00000086;
power_data[3942] = 32'h00000086;
power_data[3943] = 32'h00000086;
power_data[3944] = 32'h00000086;
power_data[3945] = 32'h00000086;
power_data[3946] = 32'h00000086;
power_data[3947] = 32'h00000086;
power_data[3948] = 32'h00000086;
power_data[3949] = 32'h00000086;
power_data[3950] = 32'h00000086;
power_data[3951] = 32'h00000086;
power_data[3952] = 32'h00000086;
power_data[3953] = 32'h00000086;
power_data[3954] = 32'h00000086;
power_data[3955] = 32'h00000086;
power_data[3956] = 32'h00000086;
power_data[3957] = 32'h00000086;
power_data[3958] = 32'h00000086;
power_data[3959] = 32'h00000086;
power_data[3960] = 32'h00000086;
power_data[3961] = 32'h00000086;
power_data[3962] = 32'h00000086;
power_data[3963] = 32'h00000086;
power_data[3964] = 32'h00000086;
power_data[3965] = 32'h00000086;
power_data[3966] = 32'h00000086;
power_data[3967] = 32'h00000086;
power_data[3968] = 32'h00000086;
power_data[3969] = 32'h00000086;
power_data[3970] = 32'h00000086;
power_data[3971] = 32'h00000086;
power_data[3972] = 32'h00000086;
power_data[3973] = 32'h00000086;
power_data[3974] = 32'h00000086;
power_data[3975] = 32'h00000086;
power_data[3976] = 32'h00000086;
power_data[3977] = 32'h00000086;
power_data[3978] = 32'h00000086;
power_data[3979] = 32'h00000086;
power_data[3980] = 32'h00000086;
power_data[3981] = 32'h00000086;
power_data[3982] = 32'h00000086;
power_data[3983] = 32'h00000086;
power_data[3984] = 32'h00000086;
power_data[3985] = 32'h00000086;
power_data[3986] = 32'h00000086;
power_data[3987] = 32'h00000086;
power_data[3988] = 32'h00000086;
power_data[3989] = 32'h00000086;
power_data[3990] = 32'h00000086;
power_data[3991] = 32'h00000086;
power_data[3992] = 32'h00000086;
power_data[3993] = 32'h00000086;
power_data[3994] = 32'h00000086;
power_data[3995] = 32'h00000086;
power_data[3996] = 32'h00000086;
power_data[3997] = 32'h00000086;
power_data[3998] = 32'h00000086;
power_data[3999] = 32'h00000086;
power_data[4000] = 32'h00000086;
power_data[4001] = 32'h00000086;
power_data[4002] = 32'h00000086;
power_data[4003] = 32'h00000086;
power_data[4004] = 32'h00000086;
power_data[4005] = 32'h00000086;
power_data[4006] = 32'h00000086;
power_data[4007] = 32'h00000086;
power_data[4008] = 32'h00000086;
power_data[4009] = 32'h00000086;
power_data[4010] = 32'h00000086;
power_data[4011] = 32'h00000086;
power_data[4012] = 32'h00000086;
power_data[4013] = 32'h00000086;
power_data[4014] = 32'h00000086;
power_data[4015] = 32'h00000086;
power_data[4016] = 32'h00000086;
power_data[4017] = 32'h00000086;
power_data[4018] = 32'h00000086;
power_data[4019] = 32'h00000086;
power_data[4020] = 32'h00000086;
power_data[4021] = 32'h00000086;
power_data[4022] = 32'h00000086;
power_data[4023] = 32'h00000086;
power_data[4024] = 32'h00000086;
power_data[4025] = 32'h00000086;
power_data[4026] = 32'h00000086;
power_data[4027] = 32'h00000086;
power_data[4028] = 32'h00000086;
power_data[4029] = 32'h00000086;
power_data[4030] = 32'h00000086;
power_data[4031] = 32'h00000086;
power_data[4032] = 32'h00000086;
power_data[4033] = 32'h00000086;
power_data[4034] = 32'h00000086;
power_data[4035] = 32'h00000086;
power_data[4036] = 32'h00000086;
power_data[4037] = 32'h00000086;
power_data[4038] = 32'h00000086;
power_data[4039] = 32'h00000086;
power_data[4040] = 32'h00000086;
power_data[4041] = 32'h00000086;
power_data[4042] = 32'h00000086;
power_data[4043] = 32'h00000086;
power_data[4044] = 32'h00000086;
power_data[4045] = 32'h00000086;
power_data[4046] = 32'h00000086;
power_data[4047] = 32'h00000086;
power_data[4048] = 32'h00000086;
power_data[4049] = 32'h00000086;
power_data[4050] = 32'h00000086;
power_data[4051] = 32'h00000086;
power_data[4052] = 32'h00000086;
power_data[4053] = 32'h00000086;
power_data[4054] = 32'h00000086;
power_data[4055] = 32'h00000086;
power_data[4056] = 32'h00000086;
power_data[4057] = 32'h00000086;
power_data[4058] = 32'h00000086;
power_data[4059] = 32'h00000086;
power_data[4060] = 32'h00000086;
power_data[4061] = 32'h00000086;
power_data[4062] = 32'h00000086;
power_data[4063] = 32'h00000086;
power_data[4064] = 32'h00000086;
power_data[4065] = 32'h00000086;
power_data[4066] = 32'h00000086;
power_data[4067] = 32'h00000086;
power_data[4068] = 32'h00000086;
power_data[4069] = 32'h00000086;
power_data[4070] = 32'h00000086;
power_data[4071] = 32'h00000086;
power_data[4072] = 32'h00000086;
power_data[4073] = 32'h00000086;
power_data[4074] = 32'h00000086;
power_data[4075] = 32'h00000086;
power_data[4076] = 32'h00000086;
power_data[4077] = 32'h00000086;
power_data[4078] = 32'h00000086;
power_data[4079] = 32'h00000086;
power_data[4080] = 32'h00000086;
power_data[4081] = 32'h00000086;
power_data[4082] = 32'h00000086;
power_data[4083] = 32'h00000086;
power_data[4084] = 32'h00000086;
power_data[4085] = 32'h00000086;
power_data[4086] = 32'h00000086;
power_data[4087] = 32'h00000086;
power_data[4088] = 32'h00000086;
power_data[4089] = 32'h00000086;
power_data[4090] = 32'h00000086;
power_data[4091] = 32'h00000086;
power_data[4092] = 32'h00000086;
power_data[4093] = 32'h00000086;
power_data[4094] = 32'h00000086;
power_data[4095] = 32'h00000086;
power_data[4096] = 32'h00000086;
power_data[4097] = 32'h00000086;
power_data[4098] = 32'h00000086;
power_data[4099] = 32'h00000086;
power_data[4100] = 32'h00000086;
power_data[4101] = 32'h00000086;
power_data[4102] = 32'h00000086;
power_data[4103] = 32'h00000086;
power_data[4104] = 32'h00000086;
power_data[4105] = 32'h00000086;
power_data[4106] = 32'h00000086;
power_data[4107] = 32'h00000086;
power_data[4108] = 32'h00000086;
power_data[4109] = 32'h00000086;
power_data[4110] = 32'h00000086;
power_data[4111] = 32'h00000086;
power_data[4112] = 32'h00000086;
power_data[4113] = 32'h00000086;
power_data[4114] = 32'h00000086;
power_data[4115] = 32'h00000086;
power_data[4116] = 32'h00000086;
power_data[4117] = 32'h00000086;
power_data[4118] = 32'h00000086;
power_data[4119] = 32'h00000086;
power_data[4120] = 32'h00000086;
power_data[4121] = 32'h00000086;
power_data[4122] = 32'h00000086;
power_data[4123] = 32'h00000086;
power_data[4124] = 32'h00000086;
power_data[4125] = 32'h00000086;
power_data[4126] = 32'h00000086;
power_data[4127] = 32'h00000086;
power_data[4128] = 32'h00000086;
power_data[4129] = 32'h00000086;
power_data[4130] = 32'h00000086;
power_data[4131] = 32'h00000086;
power_data[4132] = 32'h00000086;
power_data[4133] = 32'h00000086;
power_data[4134] = 32'h00000086;
power_data[4135] = 32'h00000086;
power_data[4136] = 32'h00000086;
power_data[4137] = 32'h00000086;
power_data[4138] = 32'h00000086;
power_data[4139] = 32'h00000086;
power_data[4140] = 32'h00000086;
power_data[4141] = 32'h00000086;
power_data[4142] = 32'h00000086;
power_data[4143] = 32'h00000086;
power_data[4144] = 32'h00000086;
power_data[4145] = 32'h00000086;
power_data[4146] = 32'h00000086;
power_data[4147] = 32'h00000086;
power_data[4148] = 32'h00000086;
power_data[4149] = 32'h00000086;
power_data[4150] = 32'h00000086;
power_data[4151] = 32'h00000086;
power_data[4152] = 32'h00000086;
power_data[4153] = 32'h00000086;
power_data[4154] = 32'h00000086;
power_data[4155] = 32'h00000086;
power_data[4156] = 32'h00000086;
power_data[4157] = 32'h00000086;
power_data[4158] = 32'h00000086;
power_data[4159] = 32'h00000086;
power_data[4160] = 32'h00000086;
power_data[4161] = 32'h00000086;
power_data[4162] = 32'h00000086;
power_data[4163] = 32'h00000086;
power_data[4164] = 32'h00000086;
power_data[4165] = 32'h00000086;
power_data[4166] = 32'h00000086;
power_data[4167] = 32'h00000086;
power_data[4168] = 32'h00000086;
power_data[4169] = 32'h00000086;
power_data[4170] = 32'h00000086;
power_data[4171] = 32'h00000086;
power_data[4172] = 32'h00000086;
power_data[4173] = 32'h00000086;
power_data[4174] = 32'h00000086;
power_data[4175] = 32'h00000086;
power_data[4176] = 32'h00000086;
power_data[4177] = 32'h00000086;
power_data[4178] = 32'h00000086;
power_data[4179] = 32'h00000086;
power_data[4180] = 32'h00000086;
power_data[4181] = 32'h00000086;
power_data[4182] = 32'h00000086;
power_data[4183] = 32'h00000086;
power_data[4184] = 32'h00000086;
power_data[4185] = 32'h00000086;
power_data[4186] = 32'h00000086;
power_data[4187] = 32'h00000086;
power_data[4188] = 32'h00000086;
power_data[4189] = 32'h00000086;
power_data[4190] = 32'h00000086;
power_data[4191] = 32'h00000086;
power_data[4192] = 32'h00000086;
power_data[4193] = 32'h00000086;
power_data[4194] = 32'h00000086;
power_data[4195] = 32'h00000086;
power_data[4196] = 32'h00000086;
power_data[4197] = 32'h00000086;
power_data[4198] = 32'h00000086;
power_data[4199] = 32'h00000086;
power_data[4200] = 32'h00000086;
power_data[4201] = 32'h00000086;
power_data[4202] = 32'h00000086;
power_data[4203] = 32'h00000086;
power_data[4204] = 32'h00000086;
power_data[4205] = 32'h00000086;
power_data[4206] = 32'h00000086;
power_data[4207] = 32'h00000086;
power_data[4208] = 32'h00000086;
power_data[4209] = 32'h00000086;
power_data[4210] = 32'h00000086;
power_data[4211] = 32'h00000086;
power_data[4212] = 32'h00000086;
power_data[4213] = 32'h00000086;
power_data[4214] = 32'h00000086;
power_data[4215] = 32'h00000086;
power_data[4216] = 32'h00000086;
power_data[4217] = 32'h00000086;
power_data[4218] = 32'h00000086;
power_data[4219] = 32'h00000086;
power_data[4220] = 32'h00000086;
power_data[4221] = 32'h00000086;
power_data[4222] = 32'h00000086;
power_data[4223] = 32'h00000086;
power_data[4224] = 32'h00000086;
power_data[4225] = 32'h00000086;
power_data[4226] = 32'h00000086;
power_data[4227] = 32'h00000086;
power_data[4228] = 32'h00000086;
power_data[4229] = 32'h00000086;
power_data[4230] = 32'h00000086;
power_data[4231] = 32'h00000086;
power_data[4232] = 32'h00000086;
power_data[4233] = 32'h00000086;
power_data[4234] = 32'h00000086;
power_data[4235] = 32'h00000086;
power_data[4236] = 32'h00000086;
power_data[4237] = 32'h00000086;
power_data[4238] = 32'h00000086;
power_data[4239] = 32'h00000086;
power_data[4240] = 32'h00000086;
power_data[4241] = 32'h00000086;
power_data[4242] = 32'h00000086;
power_data[4243] = 32'h00000086;
power_data[4244] = 32'h00000086;
power_data[4245] = 32'h00000086;
power_data[4246] = 32'h00000086;
power_data[4247] = 32'h00000086;
power_data[4248] = 32'h00000086;
power_data[4249] = 32'h00000086;
power_data[4250] = 32'h00000086;
power_data[4251] = 32'h00000082;
power_data[4252] = 32'h00000069;
power_data[4253] = 32'h00000069;
power_data[4254] = 32'h00000069;
power_data[4255] = 32'h00000069;
power_data[4256] = 32'h00000069;
power_data[4257] = 32'h00000069;
power_data[4258] = 32'h00000069;
power_data[4259] = 32'h00000069;
power_data[4260] = 32'h00000069;
power_data[4261] = 32'h00000069;
power_data[4262] = 32'h00000069;
power_data[4263] = 32'h00000069;
power_data[4264] = 32'h00000069;
power_data[4265] = 32'h00000069;
power_data[4266] = 32'h00000069;
power_data[4267] = 32'h00000069;
power_data[4268] = 32'h00000069;
power_data[4269] = 32'h00000069;
power_data[4270] = 32'h00000069;
power_data[4271] = 32'h00000069;
power_data[4272] = 32'h00000069;
power_data[4273] = 32'h00000069;
power_data[4274] = 32'h00000069;
power_data[4275] = 32'h00000069;
power_data[4276] = 32'h00000069;
power_data[4277] = 32'h00000069;
power_data[4278] = 32'h00000069;
power_data[4279] = 32'h00000069;
power_data[4280] = 32'h00000069;
power_data[4281] = 32'h00000069;
power_data[4282] = 32'h00000069;
power_data[4283] = 32'h00000069;
power_data[4284] = 32'h00000069;
power_data[4285] = 32'h00000069;
power_data[4286] = 32'h00000069;
power_data[4287] = 32'h00000069;
power_data[4288] = 32'h00000069;
power_data[4289] = 32'h00000069;
power_data[4290] = 32'h00000069;
power_data[4291] = 32'h00000069;
power_data[4292] = 32'h00000069;
power_data[4293] = 32'h00000069;
power_data[4294] = 32'h00000069;
power_data[4295] = 32'h00000069;
power_data[4296] = 32'h00000069;
power_data[4297] = 32'h00000069;
power_data[4298] = 32'h00000069;
power_data[4299] = 32'h00000069;
power_data[4300] = 32'h00000069;
power_data[4301] = 32'h00000069;
power_data[4302] = 32'h00000069;
power_data[4303] = 32'h00000069;
power_data[4304] = 32'h00000069;
power_data[4305] = 32'h00000069;
power_data[4306] = 32'h00000069;
power_data[4307] = 32'h00000069;
power_data[4308] = 32'h00000069;
power_data[4309] = 32'h00000069;
power_data[4310] = 32'h00000069;
power_data[4311] = 32'h00000069;
power_data[4312] = 32'h00000069;
power_data[4313] = 32'h00000069;
power_data[4314] = 32'h00000069;
power_data[4315] = 32'h00000069;
power_data[4316] = 32'h00000069;
power_data[4317] = 32'h00000069;
power_data[4318] = 32'h00000069;
power_data[4319] = 32'h00000069;
power_data[4320] = 32'h00000069;
power_data[4321] = 32'h00000069;
power_data[4322] = 32'h0000077d;
power_data[4323] = 32'h00000942;
power_data[4324] = 32'h00000942;
power_data[4325] = 32'h00000942;
power_data[4326] = 32'h00000942;
power_data[4327] = 32'h00000942;
power_data[4328] = 32'h00000942;
power_data[4329] = 32'h00000942;
power_data[4330] = 32'h00000942;
power_data[4331] = 32'h00000942;
power_data[4332] = 32'h00000942;
power_data[4333] = 32'h00000942;
power_data[4334] = 32'h00000942;
power_data[4335] = 32'h00000942;
power_data[4336] = 32'h00000942;
power_data[4337] = 32'h00000942;
power_data[4338] = 32'h00000942;
power_data[4339] = 32'h00000942;
power_data[4340] = 32'h00000942;
power_data[4341] = 32'h00000942;
power_data[4342] = 32'h00000942;
power_data[4343] = 32'h00000942;
power_data[4344] = 32'h00000942;
power_data[4345] = 32'h00000942;
power_data[4346] = 32'h00000942;
power_data[4347] = 32'h00000942;
power_data[4348] = 32'h00000942;
power_data[4349] = 32'h00000942;
power_data[4350] = 32'h00000942;
power_data[4351] = 32'h00000232;
power_data[4352] = 32'h00000232;
power_data[4353] = 32'h00000232;
power_data[4354] = 32'h00000232;
power_data[4355] = 32'h00000232;
power_data[4356] = 32'h00000232;
power_data[4357] = 32'h00000232;
power_data[4358] = 32'h00000232;
power_data[4359] = 32'h00000232;
power_data[4360] = 32'h00000232;
power_data[4361] = 32'h00000232;
power_data[4362] = 32'h00000232;
power_data[4363] = 32'h00000232;
power_data[4364] = 32'h00000232;
power_data[4365] = 32'h00000232;
power_data[4366] = 32'h00000232;
power_data[4367] = 32'h00000232;
power_data[4368] = 32'h00000232;
power_data[4369] = 32'h00000232;
power_data[4370] = 32'h00000232;
power_data[4371] = 32'h00000232;
power_data[4372] = 32'h00000232;
power_data[4373] = 32'h00000232;
power_data[4374] = 32'h00000232;
power_data[4375] = 32'h00000232;
power_data[4376] = 32'h00000232;
power_data[4377] = 32'h00000232;
power_data[4378] = 32'h00000232;
power_data[4379] = 32'h00000232;
power_data[4380] = 32'h00000232;
power_data[4381] = 32'h00000232;
power_data[4382] = 32'h00000232;
power_data[4383] = 32'h00000232;
power_data[4384] = 32'h00000232;
power_data[4385] = 32'h00000232;
power_data[4386] = 32'h00000232;
power_data[4387] = 32'h00000232;
power_data[4388] = 32'h00000232;
power_data[4389] = 32'h00000232;
power_data[4390] = 32'h00000232;
power_data[4391] = 32'h00000232;
power_data[4392] = 32'h000013d3;
power_data[4393] = 32'h00002e41;
power_data[4394] = 32'h00002e41;
power_data[4395] = 32'h00002e41;
power_data[4396] = 32'h00002e41;
power_data[4397] = 32'h00002e41;
power_data[4398] = 32'h00002e41;
power_data[4399] = 32'h00002e41;
power_data[4400] = 32'h00002e41;
power_data[4401] = 32'h00002e41;
power_data[4402] = 32'h00002e41;
power_data[4403] = 32'h00002e41;
power_data[4404] = 32'h00002e41;
power_data[4405] = 32'h00002e41;
power_data[4406] = 32'h00002e41;
power_data[4407] = 32'h00002e41;
power_data[4408] = 32'h00002e41;
power_data[4409] = 32'h00002e41;
power_data[4410] = 32'h00002e41;
power_data[4411] = 32'h00002e41;
power_data[4412] = 32'h00002e41;
power_data[4413] = 32'h00002e41;
power_data[4414] = 32'h00002e41;
power_data[4415] = 32'h00002e41;
power_data[4416] = 32'h00002e41;
power_data[4417] = 32'h00002e41;
power_data[4418] = 32'h00002e41;
power_data[4419] = 32'h00002e41;
power_data[4420] = 32'h00002e41;
power_data[4421] = 32'h00002e41;
power_data[4422] = 32'h00002e41;
power_data[4423] = 32'h00002e41;
power_data[4424] = 32'h00002e41;
power_data[4425] = 32'h00002e41;
power_data[4426] = 32'h00002e41;
power_data[4427] = 32'h00002e41;
power_data[4428] = 32'h00002e41;
power_data[4429] = 32'h00002e41;
power_data[4430] = 32'h00002e41;
power_data[4431] = 32'h00002e41;
power_data[4432] = 32'h00002e41;
power_data[4433] = 32'h00002e41;
power_data[4434] = 32'h00002e41;
power_data[4435] = 32'h00002e41;
power_data[4436] = 32'h00002e41;
power_data[4437] = 32'h00002e41;
power_data[4438] = 32'h00002e41;
power_data[4439] = 32'h00002e41;
power_data[4440] = 32'h00002e41;
power_data[4441] = 32'h00002e41;
power_data[4442] = 32'h00002e41;
power_data[4443] = 32'h00002e41;
power_data[4444] = 32'h00002e41;
power_data[4445] = 32'h00002e41;
power_data[4446] = 32'h00002e41;
power_data[4447] = 32'h00002e41;
power_data[4448] = 32'h00002e41;
power_data[4449] = 32'h00002e41;
power_data[4450] = 32'h000009ab;
power_data[4451] = 32'h00000086;
power_data[4452] = 32'h00000086;
power_data[4453] = 32'h00000086;
power_data[4454] = 32'h00000086;
power_data[4455] = 32'h00000086;
power_data[4456] = 32'h00000086;
power_data[4457] = 32'h00000086;
power_data[4458] = 32'h00000086;
power_data[4459] = 32'h00000086;
power_data[4460] = 32'h00000086;
power_data[4461] = 32'h00000086;
power_data[4462] = 32'h00000086;
power_data[4463] = 32'h00000086;
power_data[4464] = 32'h00000086;
power_data[4465] = 32'h00000086;
power_data[4466] = 32'h00000086;
power_data[4467] = 32'h00000086;
power_data[4468] = 32'h00000086;
power_data[4469] = 32'h00000086;
power_data[4470] = 32'h00000086;
power_data[4471] = 32'h00000086;
power_data[4472] = 32'h00000086;
power_data[4473] = 32'h00000086;
power_data[4474] = 32'h00000086;
power_data[4475] = 32'h00000086;
power_data[4476] = 32'h00000086;
power_data[4477] = 32'h00000086;
power_data[4478] = 32'h00000086;
power_data[4479] = 32'h00000086;
power_data[4480] = 32'h00000086;
power_data[4481] = 32'h00000086;
power_data[4482] = 32'h00000086;
power_data[4483] = 32'h00000086;
power_data[4484] = 32'h00000086;
power_data[4485] = 32'h00000086;
power_data[4486] = 32'h00000086;
power_data[4487] = 32'h00000086;
power_data[4488] = 32'h00000086;
power_data[4489] = 32'h00000086;
power_data[4490] = 32'h00000086;
power_data[4491] = 32'h00000086;
power_data[4492] = 32'h00000086;
power_data[4493] = 32'h00000086;
power_data[4494] = 32'h00000086;
power_data[4495] = 32'h00000086;
power_data[4496] = 32'h00000086;
power_data[4497] = 32'h00000086;
power_data[4498] = 32'h00000086;
power_data[4499] = 32'h00000086;
power_data[4500] = 32'h00000086;
power_data[4501] = 32'h00000086;
power_data[4502] = 32'h00000086;
power_data[4503] = 32'h00000086;
power_data[4504] = 32'h00000086;
power_data[4505] = 32'h00000086;
power_data[4506] = 32'h00000086;
power_data[4507] = 32'h00000086;
power_data[4508] = 32'h00000086;
power_data[4509] = 32'h00000086;
power_data[4510] = 32'h00000086;
power_data[4511] = 32'h00000086;
power_data[4512] = 32'h00000086;
power_data[4513] = 32'h00000086;
power_data[4514] = 32'h00000086;
power_data[4515] = 32'h00000086;
power_data[4516] = 32'h00000086;
power_data[4517] = 32'h00000086;
power_data[4518] = 32'h00000086;
power_data[4519] = 32'h00000086;
power_data[4520] = 32'h00000086;
power_data[4521] = 32'h00000086;
power_data[4522] = 32'h00000086;
power_data[4523] = 32'h00000086;
power_data[4524] = 32'h00000086;
power_data[4525] = 32'h00000086;
power_data[4526] = 32'h00000086;
power_data[4527] = 32'h00000086;
power_data[4528] = 32'h00000086;
power_data[4529] = 32'h00000086;
power_data[4530] = 32'h00000086;
power_data[4531] = 32'h00000086;
power_data[4532] = 32'h00000086;
power_data[4533] = 32'h00000086;
power_data[4534] = 32'h00000086;
power_data[4535] = 32'h00000086;
power_data[4536] = 32'h00000086;
power_data[4537] = 32'h00000086;
power_data[4538] = 32'h00000086;
power_data[4539] = 32'h00000086;
power_data[4540] = 32'h00000086;
power_data[4541] = 32'h00000086;
power_data[4542] = 32'h00000086;
power_data[4543] = 32'h00000086;
power_data[4544] = 32'h00000086;
power_data[4545] = 32'h00000086;
power_data[4546] = 32'h00000086;
power_data[4547] = 32'h00000086;
power_data[4548] = 32'h00000086;
power_data[4549] = 32'h00000086;
power_data[4550] = 32'h00000086;
power_data[4551] = 32'h00000086;
power_data[4552] = 32'h00000086;
power_data[4553] = 32'h00000086;
power_data[4554] = 32'h00000086;
power_data[4555] = 32'h00000086;
power_data[4556] = 32'h00000086;
power_data[4557] = 32'h00000086;
power_data[4558] = 32'h00000086;
power_data[4559] = 32'h00000086;
power_data[4560] = 32'h00000086;
power_data[4561] = 32'h00000086;
power_data[4562] = 32'h00000086;
power_data[4563] = 32'h00000086;
power_data[4564] = 32'h00000086;
power_data[4565] = 32'h00000086;
power_data[4566] = 32'h00000086;
power_data[4567] = 32'h00000086;
power_data[4568] = 32'h00000086;
power_data[4569] = 32'h00000086;
power_data[4570] = 32'h00000086;
power_data[4571] = 32'h00000086;
power_data[4572] = 32'h00000086;
power_data[4573] = 32'h00000086;
power_data[4574] = 32'h00000086;
power_data[4575] = 32'h00000086;
power_data[4576] = 32'h00000086;
power_data[4577] = 32'h00000086;
power_data[4578] = 32'h00000086;
power_data[4579] = 32'h00000086;
power_data[4580] = 32'h00000086;
power_data[4581] = 32'h00000086;
power_data[4582] = 32'h00000086;
power_data[4583] = 32'h00000086;
power_data[4584] = 32'h00000086;
power_data[4585] = 32'h00000086;
power_data[4586] = 32'h00000086;
power_data[4587] = 32'h00000086;
power_data[4588] = 32'h00000086;
power_data[4589] = 32'h00000086;
power_data[4590] = 32'h00000086;
power_data[4591] = 32'h00000086;
power_data[4592] = 32'h00000086;
power_data[4593] = 32'h00000086;
power_data[4594] = 32'h00000086;
power_data[4595] = 32'h00000086;
power_data[4596] = 32'h00000086;
power_data[4597] = 32'h00000086;
power_data[4598] = 32'h00000086;
power_data[4599] = 32'h00000086;
power_data[4600] = 32'h00000086;
power_data[4601] = 32'h00000086;
power_data[4602] = 32'h00000086;
power_data[4603] = 32'h00000086;
power_data[4604] = 32'h00000086;
power_data[4605] = 32'h00000086;
power_data[4606] = 32'h00000086;
power_data[4607] = 32'h00000086;
power_data[4608] = 32'h00000086;
power_data[4609] = 32'h00000086;
power_data[4610] = 32'h00000086;
power_data[4611] = 32'h00000086;
power_data[4612] = 32'h00000086;
power_data[4613] = 32'h00000086;
power_data[4614] = 32'h00000086;
power_data[4615] = 32'h00000086;
power_data[4616] = 32'h00000086;
power_data[4617] = 32'h00000086;
power_data[4618] = 32'h00000086;
power_data[4619] = 32'h00000086;
power_data[4620] = 32'h00000086;
power_data[4621] = 32'h00000086;
power_data[4622] = 32'h00000086;
power_data[4623] = 32'h00000086;
power_data[4624] = 32'h00000086;
power_data[4625] = 32'h00000086;
power_data[4626] = 32'h00000086;
power_data[4627] = 32'h00000086;
power_data[4628] = 32'h00000086;
power_data[4629] = 32'h00000086;
power_data[4630] = 32'h00000086;
power_data[4631] = 32'h00000086;
power_data[4632] = 32'h00000086;
power_data[4633] = 32'h00000086;
power_data[4634] = 32'h00000086;
power_data[4635] = 32'h00000086;
power_data[4636] = 32'h00000086;
power_data[4637] = 32'h00000086;
power_data[4638] = 32'h00000086;
power_data[4639] = 32'h00000086;
power_data[4640] = 32'h00000086;
power_data[4641] = 32'h00000086;
power_data[4642] = 32'h00000086;
power_data[4643] = 32'h00000086;
power_data[4644] = 32'h00000086;
power_data[4645] = 32'h00000086;
power_data[4646] = 32'h00000086;
power_data[4647] = 32'h00000086;
power_data[4648] = 32'h00000086;
power_data[4649] = 32'h00000086;
power_data[4650] = 32'h00000086;
power_data[4651] = 32'h00000086;
power_data[4652] = 32'h00000086;
power_data[4653] = 32'h00000086;
power_data[4654] = 32'h00000086;
power_data[4655] = 32'h00000086;
power_data[4656] = 32'h00000086;
power_data[4657] = 32'h00000086;
power_data[4658] = 32'h00000086;
power_data[4659] = 32'h00000086;
power_data[4660] = 32'h00000086;
power_data[4661] = 32'h00000086;
power_data[4662] = 32'h00000086;
power_data[4663] = 32'h00000086;
power_data[4664] = 32'h00000086;
power_data[4665] = 32'h00000086;
power_data[4666] = 32'h00000086;
power_data[4667] = 32'h00000086;
power_data[4668] = 32'h00000086;
power_data[4669] = 32'h00000086;
power_data[4670] = 32'h00000086;
power_data[4671] = 32'h00000086;
power_data[4672] = 32'h00000086;
power_data[4673] = 32'h00000086;
power_data[4674] = 32'h00000086;
power_data[4675] = 32'h00000086;
power_data[4676] = 32'h00000086;
power_data[4677] = 32'h00000086;
power_data[4678] = 32'h00000086;
power_data[4679] = 32'h00000086;
power_data[4680] = 32'h00000086;
power_data[4681] = 32'h00000086;
power_data[4682] = 32'h00000086;
power_data[4683] = 32'h00000086;
power_data[4684] = 32'h00000086;
power_data[4685] = 32'h00000086;
power_data[4686] = 32'h00000086;
power_data[4687] = 32'h00000086;
power_data[4688] = 32'h00000086;
power_data[4689] = 32'h00000086;
power_data[4690] = 32'h00000086;
power_data[4691] = 32'h00000086;
power_data[4692] = 32'h00000086;
power_data[4693] = 32'h00000086;
power_data[4694] = 32'h00000086;
power_data[4695] = 32'h00000086;
power_data[4696] = 32'h00000086;
power_data[4697] = 32'h00000086;
power_data[4698] = 32'h00000086;
power_data[4699] = 32'h00000086;
power_data[4700] = 32'h00000086;
power_data[4701] = 32'h00000086;
power_data[4702] = 32'h00000086;
power_data[4703] = 32'h00000086;
power_data[4704] = 32'h00000086;
power_data[4705] = 32'h00000086;
power_data[4706] = 32'h00000086;
power_data[4707] = 32'h00000086;
power_data[4708] = 32'h00000086;
power_data[4709] = 32'h00000086;
power_data[4710] = 32'h00000086;
power_data[4711] = 32'h00000086;
power_data[4712] = 32'h00000086;
power_data[4713] = 32'h00000086;
power_data[4714] = 32'h00000086;
power_data[4715] = 32'h00000086;
power_data[4716] = 32'h00000086;
power_data[4717] = 32'h00000086;
power_data[4718] = 32'h00000086;
power_data[4719] = 32'h00000086;
power_data[4720] = 32'h00000086;
power_data[4721] = 32'h00000086;
power_data[4722] = 32'h00000086;
power_data[4723] = 32'h00000086;
power_data[4724] = 32'h00000086;
power_data[4725] = 32'h00000086;
power_data[4726] = 32'h00000086;
power_data[4727] = 32'h00000086;
power_data[4728] = 32'h00000086;
power_data[4729] = 32'h00000086;
power_data[4730] = 32'h00000086;
power_data[4731] = 32'h00000086;
power_data[4732] = 32'h00000086;
power_data[4733] = 32'h00000086;
power_data[4734] = 32'h00000086;
power_data[4735] = 32'h00000086;
power_data[4736] = 32'h00000086;
power_data[4737] = 32'h00000086;
power_data[4738] = 32'h00000086;
power_data[4739] = 32'h00000086;
power_data[4740] = 32'h00000086;
power_data[4741] = 32'h00000086;
power_data[4742] = 32'h00000086;
power_data[4743] = 32'h00000086;
power_data[4744] = 32'h00000086;
power_data[4745] = 32'h00000086;
power_data[4746] = 32'h00000086;
power_data[4747] = 32'h00000086;
power_data[4748] = 32'h00000086;
power_data[4749] = 32'h00000086;
power_data[4750] = 32'h00000086;
power_data[4751] = 32'h00000086;
power_data[4752] = 32'h00000086;
power_data[4753] = 32'h00000086;
power_data[4754] = 32'h00000086;
power_data[4755] = 32'h00000086;
power_data[4756] = 32'h00000086;
power_data[4757] = 32'h00000086;
power_data[4758] = 32'h00000086;
power_data[4759] = 32'h00000086;
power_data[4760] = 32'h00000086;
power_data[4761] = 32'h00000086;
power_data[4762] = 32'h00000086;
power_data[4763] = 32'h00000082;
power_data[4764] = 32'h00000069;
power_data[4765] = 32'h00000069;
power_data[4766] = 32'h00000069;
power_data[4767] = 32'h00000069;
power_data[4768] = 32'h00000069;
power_data[4769] = 32'h00000069;
power_data[4770] = 32'h00000069;
power_data[4771] = 32'h00000069;
power_data[4772] = 32'h00000069;
power_data[4773] = 32'h00000069;
power_data[4774] = 32'h00000069;
power_data[4775] = 32'h00000069;
power_data[4776] = 32'h00000069;
power_data[4777] = 32'h00000069;
power_data[4778] = 32'h00000069;
power_data[4779] = 32'h00000069;
power_data[4780] = 32'h00000069;
power_data[4781] = 32'h00000069;
power_data[4782] = 32'h00000069;
power_data[4783] = 32'h00000069;
power_data[4784] = 32'h00000069;
power_data[4785] = 32'h00000069;
power_data[4786] = 32'h00000069;
power_data[4787] = 32'h00000069;
power_data[4788] = 32'h00000069;
power_data[4789] = 32'h00000069;
power_data[4790] = 32'h00000069;
power_data[4791] = 32'h00000069;
power_data[4792] = 32'h00000069;
power_data[4793] = 32'h00000069;
power_data[4794] = 32'h00000069;
power_data[4795] = 32'h00000069;
power_data[4796] = 32'h00000069;
power_data[4797] = 32'h00000069;
power_data[4798] = 32'h00000069;
power_data[4799] = 32'h00000069;
power_data[4800] = 32'h00000069;
power_data[4801] = 32'h00000069;
power_data[4802] = 32'h00000069;
power_data[4803] = 32'h00000069;
power_data[4804] = 32'h00000069;
power_data[4805] = 32'h00000069;
power_data[4806] = 32'h00000069;
power_data[4807] = 32'h00000069;
power_data[4808] = 32'h00000069;
power_data[4809] = 32'h00000069;
power_data[4810] = 32'h00000069;
power_data[4811] = 32'h00000069;
power_data[4812] = 32'h00000069;
power_data[4813] = 32'h00000069;
power_data[4814] = 32'h00000069;
power_data[4815] = 32'h00000069;
power_data[4816] = 32'h00000069;
power_data[4817] = 32'h00000069;
power_data[4818] = 32'h00000069;
power_data[4819] = 32'h00000069;
power_data[4820] = 32'h00000069;
power_data[4821] = 32'h00000069;
power_data[4822] = 32'h00000069;
power_data[4823] = 32'h00000069;
power_data[4824] = 32'h00000069;
power_data[4825] = 32'h00000069;
power_data[4826] = 32'h00000069;
power_data[4827] = 32'h00000069;
power_data[4828] = 32'h00000069;
power_data[4829] = 32'h00000069;
power_data[4830] = 32'h00000069;
power_data[4831] = 32'h00000069;
power_data[4832] = 32'h00000069;
power_data[4833] = 32'h00000069;
power_data[4834] = 32'h0000077d;
power_data[4835] = 32'h00000942;
power_data[4836] = 32'h00000942;
power_data[4837] = 32'h00000942;
power_data[4838] = 32'h00000942;
power_data[4839] = 32'h00000942;
power_data[4840] = 32'h00000942;
power_data[4841] = 32'h00000942;
power_data[4842] = 32'h00000942;
power_data[4843] = 32'h00000942;
power_data[4844] = 32'h00000942;
power_data[4845] = 32'h00000942;
power_data[4846] = 32'h00000942;
power_data[4847] = 32'h00000942;
power_data[4848] = 32'h00000942;
power_data[4849] = 32'h00000942;
power_data[4850] = 32'h00000942;
power_data[4851] = 32'h00000942;
power_data[4852] = 32'h00000942;
power_data[4853] = 32'h00000942;
power_data[4854] = 32'h00000942;
power_data[4855] = 32'h00000942;
power_data[4856] = 32'h00000942;
power_data[4857] = 32'h00000942;
power_data[4858] = 32'h00000942;
power_data[4859] = 32'h00000942;
power_data[4860] = 32'h00000942;
power_data[4861] = 32'h00000942;
power_data[4862] = 32'h00000942;
power_data[4863] = 32'h00000232;
power_data[4864] = 32'h00000232;
power_data[4865] = 32'h00000232;
power_data[4866] = 32'h00000232;
power_data[4867] = 32'h00000232;
power_data[4868] = 32'h00000232;
power_data[4869] = 32'h00000232;
power_data[4870] = 32'h00000232;
power_data[4871] = 32'h00000232;
power_data[4872] = 32'h00000232;
power_data[4873] = 32'h00000232;
power_data[4874] = 32'h00000232;
power_data[4875] = 32'h00000232;
power_data[4876] = 32'h00000232;
power_data[4877] = 32'h00000232;
power_data[4878] = 32'h00000232;
power_data[4879] = 32'h00000232;
power_data[4880] = 32'h00000232;
power_data[4881] = 32'h00000232;
power_data[4882] = 32'h00000232;
power_data[4883] = 32'h00000232;
power_data[4884] = 32'h00000232;
power_data[4885] = 32'h00000232;
power_data[4886] = 32'h00000232;
power_data[4887] = 32'h00000232;
power_data[4888] = 32'h00000232;
power_data[4889] = 32'h00000232;
power_data[4890] = 32'h00000232;
power_data[4891] = 32'h00000232;
power_data[4892] = 32'h00000232;
power_data[4893] = 32'h00000232;
power_data[4894] = 32'h00000232;
power_data[4895] = 32'h00000232;
power_data[4896] = 32'h00000232;
power_data[4897] = 32'h00000232;
power_data[4898] = 32'h00000232;
power_data[4899] = 32'h00000232;
power_data[4900] = 32'h00000232;
power_data[4901] = 32'h00000232;
power_data[4902] = 32'h00000232;
power_data[4903] = 32'h00000232;
power_data[4904] = 32'h000013d3;
power_data[4905] = 32'h00002e41;
power_data[4906] = 32'h00002e41;
power_data[4907] = 32'h00002e41;
power_data[4908] = 32'h00002e41;
power_data[4909] = 32'h00002e41;
power_data[4910] = 32'h00002e41;
power_data[4911] = 32'h00002e41;
power_data[4912] = 32'h00002e41;
power_data[4913] = 32'h00002e41;
power_data[4914] = 32'h00002e41;
power_data[4915] = 32'h00002e41;
power_data[4916] = 32'h00002e41;
power_data[4917] = 32'h00002e41;
power_data[4918] = 32'h00002e41;
power_data[4919] = 32'h00002e41;
power_data[4920] = 32'h00002e41;
power_data[4921] = 32'h00002e41;
power_data[4922] = 32'h00002e41;
power_data[4923] = 32'h00002e41;
power_data[4924] = 32'h00002e41;
power_data[4925] = 32'h00002e41;
power_data[4926] = 32'h00002e41;
power_data[4927] = 32'h00002e41;
power_data[4928] = 32'h00002e41;
power_data[4929] = 32'h00002e41;
power_data[4930] = 32'h00002e41;
power_data[4931] = 32'h00002e41;
power_data[4932] = 32'h00002e41;
power_data[4933] = 32'h00002e41;
power_data[4934] = 32'h00002e41;
power_data[4935] = 32'h00002e41;
power_data[4936] = 32'h00002e41;
power_data[4937] = 32'h00002e41;
power_data[4938] = 32'h00002e41;
power_data[4939] = 32'h00002e41;
power_data[4940] = 32'h00002e41;
power_data[4941] = 32'h00002e41;
power_data[4942] = 32'h00002e41;
power_data[4943] = 32'h00002e41;
power_data[4944] = 32'h00002e41;
power_data[4945] = 32'h00002e41;
power_data[4946] = 32'h00002e41;
power_data[4947] = 32'h00002e41;
power_data[4948] = 32'h00002e41;
power_data[4949] = 32'h00002e41;
power_data[4950] = 32'h00002e41;
power_data[4951] = 32'h00002e41;
power_data[4952] = 32'h00002e41;
power_data[4953] = 32'h00002e41;
power_data[4954] = 32'h00002e41;
power_data[4955] = 32'h00002e41;
power_data[4956] = 32'h00002e41;
power_data[4957] = 32'h00002e41;
power_data[4958] = 32'h00002e41;
power_data[4959] = 32'h00002e41;
power_data[4960] = 32'h00002e41;
power_data[4961] = 32'h00002e41;
power_data[4962] = 32'h000009ab;
power_data[4963] = 32'h00000086;
power_data[4964] = 32'h00000086;
power_data[4965] = 32'h00000086;
power_data[4966] = 32'h00000086;
power_data[4967] = 32'h00000086;
power_data[4968] = 32'h00000086;
power_data[4969] = 32'h00000086;
power_data[4970] = 32'h00000086;
power_data[4971] = 32'h00000086;
power_data[4972] = 32'h00000086;
power_data[4973] = 32'h00000086;
power_data[4974] = 32'h00000086;
power_data[4975] = 32'h00000086;
power_data[4976] = 32'h00000086;
power_data[4977] = 32'h00000086;
power_data[4978] = 32'h00000086;
power_data[4979] = 32'h00000086;
power_data[4980] = 32'h00000086;
power_data[4981] = 32'h00000086;
power_data[4982] = 32'h00000086;
power_data[4983] = 32'h00000086;
power_data[4984] = 32'h00000086;
power_data[4985] = 32'h00000086;
power_data[4986] = 32'h00000086;
power_data[4987] = 32'h00000086;
power_data[4988] = 32'h00000086;
power_data[4989] = 32'h00000086;
power_data[4990] = 32'h00000086;
power_data[4991] = 32'h00000086;
power_data[4992] = 32'h00000086;
power_data[4993] = 32'h00000086;
power_data[4994] = 32'h00000086;
power_data[4995] = 32'h00000086;
power_data[4996] = 32'h00000086;
power_data[4997] = 32'h00000086;
power_data[4998] = 32'h00000086;
power_data[4999] = 32'h00000086;
    
end

endmodule